XlxV64EB    fa00    2fb0*���s.��\�P�]�k.O�5仑q�S��I��T�>��ұ��x#Ԓ�lU�vM�����6�����1�C&�����E�?��F����:�c��\�g2�����4{Cج�����K�SG�!��r�����1�
N����>#q_X��6�ә�����hD}�W=d�_��U��s�*��Q|^��$��a�.�D'zY�0�SL!���U#_s^��N
��FɒƓ�vܻx?u�w1���W�E[���V��)c(�j?<5p�5��cnڛ���k(;��[o�4�D�]��̟��"�ڿQ�Z ���N���ЩyjH��C`QrĿ��i컅��o�E��$����'KD���Rf��𵓴-�R�8SV��4����D�=aa#�d��}�i�榆#�t�����[��)���ߓ#����ѱ93�ρi@�j�p�/�g3�
~y�m6���M`h@�p�P�n:��
�y{�*��׳���AqW1��	cU�HRos�㸠R���čJ����m�}��t>k�O��$��r^�~��2�Hi%>����Dm��A�4�"�x��UF�i�
*|��P�kIF`��n �t��m���#���D?j�bSl".n (C]O3�Q�����u
O�;&^�f�/��}s������%3�f�)��Pvy�@ӂD�?���������m��
����R,�د^0:0�Kx�e�d��ى4[� � l����l�^{���]p�I:#�#)a%z�{�ȰiR�������'� B&�mwY�l��-�Hhr��J�ؠ�4�C}��בc��
8�#���#�T�4m@z��(��kO�֮řk��&CB�8wV��w9W�1�p�?1*	R�d��4�����h�3�ɀ���8*iz��rj]��7^W��r'�k����Fv�9�\m�0t�XJ�N�%n�����$�6�b_�kF>邶��#ű@�ug�$����^��w��Rݸ����<�+��҄�V:3���1iGl�S4��/F�wϾ}�ֽ�|�U[}|O!5D*��1=��>����#���y�9X�X�I�ij�W܅�Ѥ�<���Н�`Ӗ��>Up������:̅/N9�o�8�6�������CE�h@��ޝ*b*�.�P�Yʶ6a�1�������l�Cu��� ��}� ���qH�7��?�ꭗ>׾UVd�D �ɱO�ĲM_�H,�%���U_2�1��SQ��u\,,�$]�<����1
|uD#G��櫓v�މ����LR{�&��y/ϙ��sp�q7�c)�_ot�+!-#���dN���<k��&>5�����ק����md��.���tr��ĻM�츀6��M1:O]ܮ�6#�5|l�o���,�!܉�����v@e��Ua4>�x��V� �<s�`P�&��8	��r����ˠ��7�8s�%2	"�*%d>���Z��_���H'Ž.hW\�$���s^�Uw���ĵ�/�Vj0;��U@eֽ���:��cLó�>AX�G�X��R�6�u�������ķ�i���VD��y1���O]�jb�T34ݧ��r�aݜMr�T`UA9`�7�|*s����dmj�i=����Z��*f�����h�B�<l0xr��q?$�ud�V����D��FS;@�ig�NU��2!� B��s(��~�Rn�����*8LW�7U��@|u6����\и��_D�)x��=|\H#�	��-c�U�/��'�zϢ|y���+�f���Ɏ��l�CLc?�����, 5l� Y�4�A�Y�U. ��>��pn���XA�W���9���f�B�UyW�{�D`A�_0��Y��ne��9js.�j�z�苳�kxTO*��E};p�H����B�m��V��>���׬���\�������>CZYՄ�LH���K%3���	d^%�u��-R#3��H_�N���0�v�R���,_d/g�ܶæ'8(����§[�sK��%J���Dn������'�(WiL�H�0�	���dߣb�r�sJ ��T��>E�>+�0S+���x�8��/�=�Q�Z1!���� ��q��"i�k�Z ��}R�YJl�è�ؓ���^�¶z>��ը�hQ�Yk�O��w  ��>E��m0�@���D����-w������Q���1�w'8����Ǎ&9�*\_�:g	|%����,qn�I�B�(�Z_{0���Us#Q����B��e2f�m�����'E6�� �?.'�MХ�I��s ):���R���+!]o��=j	����~`L*v���l���Ђ\N�����\����R��@ݐ���[ �6T���;o�
b��V�ڹ�|GJ�{��G�Fי��mɖ	��퍾�*ぉ���s�[�+���}�F�%����(e��?L�-�?8}��U�ǯ�ڽ(�t�j��t9�+�@KT����p3�ٺ�Z��i��Iz_�gTs����	v��rc�V���)d��p�Yl��x�����NP֒M�'�6t4^��!VYI'����\���(����ģ�L�::�d0��m�('i
L"<�������U���Ym�m!�)kXW�}�)���W�d򐐰oa��������kR���Z��(��9�EN�X��U�Qm���22����LL|{���Z�lu�k$�Q�p_h����4i�����������l��'���aU�����'sd�RZH����0���N���� ��\�����?��/��,���A�'�U��_�i�Ϥ �X�M���{tS�A\����z�h��1$�3���e��N�WeԯGf�-��n&9;���ۃ�S%��_�r�&,hh\��k��Ui'KG2�Ss�a�W0a�I)����������f�����g�e�G���5^�L�j�X2P�Y�r�9�<��
����cv��wTV����WKa��~a%P�yR?sF�{A��
���{r|�<�:���lݲߍ���B1͟#�1���3�:,����6��n�8�W�[,V%N�Ι�eC�|�!UA�B�"f2!\ᐯ��B��!�b�ӳ�i;~u�ɲ��"<H�dV�u�­�8���bɄ;�G-6J����C(�]F�T��w���/����ќ�sZ����K�Xd��h��HzJ�3k�Y���� bd��6lAH�"Y���6�����-�=��v��������������|�7�	�J��堢iBh%�f!��(�^j_������7�H�����%Ky��� R�;M�9m}���xy~x��]?�r�M��HY���߸_8���>��&ڴ[��vh��po��ܦ^�����$�����ˎ~ Fne��_TO�k��c���)�B�ɳ��&9KlE��(=�r�L>ߑV��g�9�Յ�z7�Ou|�xzl>T}Z eB҈���;f2�@���Lf���x�WD�B��;RM�%�۲��H�d�u ��yd�d!���~�lF���e����w�Bw��� ���x�|x)�3_��3
y�+|s�AwG��@�1w(5M�{e���E�R���"�[$pOyNq^|���о=��'�kJڲC�H!��\T�jJ��M2[9y�+&؅!:RMr�-n����X���;�K�WQB�g��K�L��?�)�c48/��#�<	���}=����4L���D$�3k��u��t)���=�R��"M<�ܷ`2�XOuL2̜��̪e �أh"�6n7
�LK���u����	{�z�XU~Ų64�s�}<g�
L��q^A��dȁwʍ�m��*V6D��υ�ϧ&&���Dh��`�;<q�Ǉ��mpár��AnH�sf�3]��Ba�2�!��@����n#@��Ӱug5I����a˙Ve�y�n���-�]�������[�k�X�3Ə�4��%`�q��)v�\����>����v���Ez@�P0Gmޖ�s9�{�?��9�ݯr�A���8q6.���$M�2�ҟyyL]�nNW�3:4H�I �zۍ��Z�����̳��'�h��ˡ]x�Lx'�}J��6`�@��ѻ�e���� t��XK쉖X'kz�������x�;&+D�0��;-��Ն%�B�q�����qƓ�Z[d�g���;5�~p�"��MUu�	����W"���$��Oٻ8o��{���]F3۲�Cg��aV���U���=O���Hu�g�:��!D��� x����.���{��|T�\�'�ߐ�3\����ϝ_������ˈ&��!��ۋz�̙w�O�Lx��'c��_Pgr4��`l��uzOH�(&�ɒϪ.�Ƌm�ʙh��PV��>�6sr!�� Ex���LL>�&�H����
�XpC��~ܭ�Lf�~�CfH�<:��a���+d�3.f?j�!� ��Ʉ���x�k��wA"bf���Ci�7���L��'��$ts�cfخ�ZȀ���@�>7��#.�8��/0�� p�]�Ĝo���sQ��(�0����щ�bw~�)]�)^=j0����;vSE�ټB�$�@����ꝵ`p��Wvtq|bw��0�=Z��K�p⢲��լ0*yd��[�k�F NF��y~�FCa&��ړ��rCV,�Wj�Sdi�lD�.a�����bã��Z����B��b4*뼳/�f��b������s�BQ���~�� ����""��vy�6D�.��C��t�*g��W	2�]�K:l��dl.��S� �EEg��>�4&��Q\����q�H7�֎���ȕB��?��5M?�����zR�#��c�DSc�K6�]��/���z�b*Ի�@�v"�oχ���K=�3r�w���:T������֫����[��,�sJ6�ָBK�0nU>���7�cݸn�/P����o���%�Vy��V��6xɅ����A��'�B���C�r�ɥ
�)��u"٧��-�<�7l���@.H�4��/7��[!4u��w���~�|9"�爐�����̩��r���on
j/�3�t�p/���s�m�GǮ,�P����4���������d��7A31�G$9�����A{e��l�1��hY��];G$
Ŵ	F�X]Ӕ����/�٬I+�P9T�ʎ���^^����CGUj�K�k%5C����._���->�o�>�?���W��v-=�Aɏb����n�v5�NL22s��*Nk��/�v��\iiL{߿˗���4�({8��i.c�w,}C�6L�J����}���0�-��xn�ó�/l;�A�Y�NEt���.v!RA�v!c�)لS�;�A�[���0�P�F��&b�,h�3yU���AN��{�O�I��* `;�R� b���A�X-4��izp 8M��U�,=Do�ĻE8�<QY �喤p�8���-'�h����1)«�>\V�[g��S� ^�����Lu�Oa�&����V%b|
����w65f�[�t�wXB��F � df]������Q:��;���	�.�/�<�w�BJ��q��
fS���X�,td�ø$\#Y�kCy]��_��&�H���B4��#���g��e>sd��8�;�#u��G�O��v���1��H-i	d�p#�͝�ju�F1I	�f�Л��/K��/�F%�P=�{�PZ����=j�;ޫ�W����3�A��걛�)n�p!��3H�b���4�F����ux�뼫`(�\=b���.�P@*N�>6�,���̮ϧ ��ׇ�ڪ-ܟq}ռ�)��~�F�=��3���#�_�P"�lYj��彙cs}����A�L2H�v�(��$��4�E�R�?:Gd���6w����yq�vHW#_�6S&k��R�ʙ�򨺅N6��0@������=������l/��o�V#R���Ra�P���8�2�?Ք��*�t@x<p��Z��E�*�J�F,�,�qH���{�}׹o����A;�ג�tHR��u�)��8���X�A�Y���}�E.W�7RJ�R�~�:��dH�z��g�À�l	�Y��ٍ���: #󑟲4��f�R�%F4vj㙂6Ǒ� ��k�h�r@SƽǇ��C[Wh^���C]�	�a(o�N�}�]2�x��{�G
�)e�r�����������;,��3{��kS�OQ�ҕ�w�����5�׉
y�j[$����h`����¹��^���q�E�V7�j<7gq@���j\uf��J�ٱ��}����`RN�`â�<1�
ʵFu��3����Cw5	UT�@��:�o�f��ɸ(���Q��|ZD��֘�±�3`(�]O���Bd����x��?�#נ�ʶty�$�L���jav�)0���X輤���s�u���b����,��'6��O%yܺ����[g/p"�Q
�ݝ�2�H�Ȏ
���0��6Ó&G��Sa���ݮ\��#�T��m#�FcA`=�%0�_fl��M�ի�r6�d)�`�ӵ�K��kH�l��v���~HMV%MØ'�j��&�wP�|�AC}I��We��z1]�=���P^���9#�G�Z���?�~��4�-<�j��򟽴����`��b�l;ҧc4���5R�5Ky�~D���Ĉ�¢�EkU�s�i����:x�g�jO��N�$�qJ��%^+���`5�F�b����E�9�Vfz�EE�����*:�%b���U���ts�ά����l?�ʫa[��&����������Xn�ۋ+vg��-x�#����?��������D.t�m>L6�sS�v��B�U��$�,��f��9��v��]��,]��C�N�O��sH���B����\;2�l�-XX���B"9���~wS��g�@��+[:��ՑfV�yi����4s	�J[��a�%@R�W�F�D'n���h�(�,�f7B�񰇕���*��Q=|4U(����n�B������yD~jd��z<wͮ~��^����X�,��'���V�L"~�ݟ���9�ҁ����U.Zo�L�L�� ��|��B	$�#�e4�>�m����>_5-ӐP�JA�6�Fj���iP1(�� �0��l�������	����ER#Y�$�S�ƒ�=_io�{h��=OT�j� ����V�Ő9{�7)�lf�[�����ꋋ�j��$�Y�UL���l֍������;Od�Oty���|^AP���KϗK�b�6��n<����F�}KI������ �e�5le⢂j�i��Wt���L��U�Y����^07�ga����VA����P����XC�ZN�����L�]�h9)?�c�	�ŵa�_����/A�]\��v{g��m]�Zx���G�)��lRU�]Søjs���*"�]'��E�ꛔ��|��}=���d�!7K���0xw;ˏW��E�q�>��f�*�f�o�����e������+����������z��G11�5Ɓd��7�s����5D]ћ�9���~��}7��_xKt����VE@���/��i���D��]r[���[ٜ�BM�of�����D����wh?�p٪�Z�R��2�&5�߻!�[�q�H���o6�}��)4QLD����DA����d�N��y���e	;�VrC=��)�1zK���֙}��:�F4ɑ��ET�du����w��%*���d]j�Ǟ�Q���Y��4���T�ٕT�J!l͂�,�0!'�l:Yv���N�d�!��Iu��-І��b���&�X%�(҅z��\�x��~�ς��1�c㿾79`������`�g��5$UoWH�����z�k�'(�b+��<7�x�i1�(j������8�+:g�����&�
/��&��+�q���A	��/��P2����봶������|�4�zts��`�"_�n�3���4��nt�b���]�7̃�T�W���j�YC=��|���f�`���&V��,i�\-A/��mqq��vy�&Aߗ�
Τ 	��t��.����K�G	�f���N���K�R���/@��@@ �'_��Ah�OɤX���W4Z'�cK[�u]�����Y�,�t]��t�<I��M�@���s���	�k1j�x�t"���@|{E��֪��n�B���0'O0�s��P��ʂ�Q�/��(0�Ŝ�a�Ҵ�QlUt��qn6�>�x!��N��H���r��^��U�O{V�+��L}�5'��n(���4�?�k�d�Dm��գ/���m1�ɀ�m(�����"B)E�o�h;�f�ȁ� �|�,)�u�k"C��v�CΌ��8��3ū~�'��gĽ x(��40�t����^����_>Mx�]��FOoTaW���r}nz=�Up�#Ⱦ�6�`�l��K����+�	V��,:�r~V�>�j����
���;��+fU�!k��)�Ʈ���M�c�ْ ۣ�NF�g�W�S������L�D���X{��*AG$o�.����'�T���86�iǥT�#�Q�DW��,N"܃���ڞ��l��;F�|�&�f��6��V�̞ܺ��CE��.R�~j���F���p��J����(���Q�6?�nfz>�s^��6/a:~tt�d�Z�r��m�W��`-:10vPbg��^T��_7Hr>	� ����{u1�ec*�Qc~*M/%$���'�Q;W\w�f��W2��X?9fF��Zc00��<hU؆\$��4��6�H��,߆�-����!��L�"�8�,B�CX�.^j�<�PX������D��J��t"1a�R��2��z���d�QL|����y�Gy[������){!�=��O����Ň���mI���0Ԝ*���7�aƨ8PkŨ�?7�J�;�ڵ,[���{Ss�>v�Uk�x�6@��G�"(�@I�5)��AuPu޽��Uد��o 6ɥ���6'�L�bE�#|W�@�Hz���N���-��c��D*�lJ:�t��]���e�z�����Ү2U>��Wj��/^L��om�0{�`DR�kF�V�`��/ 1��>����G�F����V#���[m�<�%��|B{aǒ�����o4X6�`5�~#�+�M:�Y�5�5��Y�bPn�tr�kW�k���zՊ�5pU�����Z�ߏ+�Wj��S�p ؉Gl�>�l>�����w`(2����w����I��Lvl��XʮLg�!1�d�n���e]�rU�w{B�'�1�Kuu��������>�z�5juɐ�4�)&���[%���9]��n���ʣ�/5��%U�����]σ%��&���gEe�k�/o��'�?;���gpf�v�yC��+��Ղ6h���;��!�٫��9� ��@�m ��}`�ax
�hW�H��[�L6묶c���qeF����59nD��O����$z��) ��lRx��O<�Z9���,ʠ4�z[��i���/�T_�����E���+c�������n7�\�����.q���u��Z��f4�bBa�?�9�p��a���߶+o/2� N~\P�bg~������_p��S׻\�d� �C?h�Q#��}��['���s*-,[��F����֖��2fTg���䂇	F�a�7&��0�M��G
��($���
ˆ-��a�8���,�r�Zj4�aր��0���t+
�B���遮��7���	��#+Y��bk����ϒ�d��F)R�S�6��v��1��U:�z�a��z:e�AAi�����(\�p��wv��V���:�'=���@�$Шc+����8Ё�ݰTXӣ��f���Y�yfG
��w��wiF��x�:=됛�p6K���%bB��%P�ab����2�slPz}7��x7z���غ��v1��"F�Do�����BKbI�ܢ75�o-.ǿԵR��Dy���%*{N��*>�rB��Q���~9�+ׅ�VR�� ���J���QH:�� Нc)����#�~3��Y�0���dOX}��!3iZx��1�$�����3��?]W���J��v����6�kK��̤X(3U�M�)���й��DX���Q�w��� ȶ���`I?�q�b�lE�½J^q��i_�pD��K�\��eN�}ȓ�@��\��+'��	D݋kK�l�!#��jh���*�RzA{���� ���Oò��d�^'���N�GI��%�_޸�58�g����]=�
��	���_�����C(���ֺ�|���|#���K5�ҋܜq�'���^2��y��`���[�^�XR�;Rb����=ξ�Q+P;���w\ll��ʪ�ɾ ��h�B�,���A��BG�q�Z�_���ou�"�%$$_��;|��4&ݮ�@!��.Q;��k0>�x��J���B1��E`�FFkl:�to"�Fao{a�dL$h�N��,��qʳ��;X1��_����B�x�|��6�ŷB�[���I��S^�6T���	�'��ٰi˰[T��߶tXo]e�-]#s���u����PJ>��3�R��e�������`*&N+���GU�� �[2�j��;���N^�� ����6
�ݔsΝ�Z(��� R��M&"�W#��Đ�a|n8ᴛ�~��	c��j���@ϼ�U���z�J��}tAIӰPBPr���ق�D{,9�۪���X�[jbWk����*Qa6�$�.}�/��c�a�)�d_���My�Rټ!+;��j:�v�Ӫc�-�"87���[����aS����إￌT�����Zͬ��	M� /����e�E�ٛ-P�m�T��lRo�\�eG�u�D�-ʊ�b3M�]�`���^�C�G��mq�@��{䒋�m��,���C��ğ,NpJ���o��&ڈ�J<����i��-������t��ˣ�d�yѮ���=�C2S���x.�� k:B�O�N�i���T�B?A�*��]��Tj��G�6EO�`����}'�Rh�F�n�"��O��c�f��NA�*p��]�]��bN'.�ό��O(��$�RLW(�jOwub�`X0�$�T+��o��࿛&���6H�`9�;jC	v�B�F��P4��U���G����$��Ǡ����-�����B��H�io��� ��#��4:�����(�Z=ʧ:��3uf�H�J��¡ow�{-�p�M�B�������4f@�Y^�޼f��؀q^KpC��;�2IoA����O&X-�+4�NbL]ȓr}�&:�6pC`��� (�?�Aء\�o�戵�HC�0U�~����T�}�aSa70+��Ln��A��Z=z$��>�,�}h��l\�`��.�Ĥ��;xi��� U`1Tug烩���o����rUn��`�e+%ƀ�S����p�}�e���,�X�e���9u��l�bX�}����ܩ_��k�~h�n:tC>�����8�R*���«�D�mN���#E���@f��=7���G����rj�r�w"eRЄ	K��l�L��RxI?I���G��q�!ri��k�7��)�����v%H��畒ݖ^���w�J��C. �%A�	[��{(mD:fl��'�"�&u�>�����~���kj�	���$9�l��Ҏ������v��N]49�>��s��,��ȇt"B��R�'�-B�cż������]�'
���A%�v���˞mQ!W�U �X��x�W�  ��aI�Xcw�J��ea�� ��wn����X�\V8?�h~Q�V��.n���3A����Mޢh��W�W��_�K�_�
UB���>=a��~�!d�x�{!q7W��ߵ��8��r�x�A�M�t�Y$�����-�8��n�A�f���V/��i���m��k6Ɲ�z]���7V+��cۊi�#�^A�c�Wg$��]�DO�[�;�.D�'��L��ُ�8e.��~��cJ�[Rx~Rn���d�иg���ܼ�%�J�S��z$�Ю~"�%�\��sK�uS�}6T���$O��L6HP*�t.:6>U�W���5v�������*Ӛ4��潚�����ߋXlxV64EB    2add     970�����@��O+yi\��:��ǿ�6�9�����|p���ˤ0G/�G"]�Ai�JT�_��g0�8�YqC=0�j�L��yMIW�=�$�#�؆���~}�ĂB�?r���W�||�b�D9(��DH^m?lN	m����?ߡcĩ?��$Ia,�1���3�ÎZ,�ؗSEd(\X��hs��de���P	O@.:�<2�̔c[i�^ze
�&р0�V�τh�O����L��[1��.�;�_��L1��sc��iv���͸�������L�A.�
%��	I2{��t���crSɬ`���b�亳
]jA�Xܩz5ܖ�W�  vao���y}U1O��b�����s��(���l�������!r�!.�o�<Ե I���*�D��̉;��p�^��j|�E�lp�^DPi�^�;�9N��G�@ Fݻ?��i�t��@��ܷx!ȿ��y�u�2ILO��]�8>�O�`��!�#�����C�D#w���U�L-���1N�h�;�R�k� f#-� �eL|�i�ߖ)��e�@�����Q���r��Fp��i�m�f�Ȕ��(�1��C�Lh��c۱%�M�/{��J�a����0�9\�B<@����}�&���ed5%ײ��ư_(�\��:��"�c�[7]-���H2����]��˂�04�
�	^ǓH��HA���t�tT�м!�ҜT��d�Ɇf�6���	_��~���� _Iv����4����bjpy��Lg��&�631'e�-񽃀ELR&�������&���e;�ǡ`�j(I��SGw� a&��/V�ߔ�Pb쩂���9��-���n��$�Y�<�����N���|YgT. ��3�QoG6��'���H��Ģ�A(� wi�����QҐ��9kq���
4�
��{	л"`Q!R ��hQ�k 6��f��G�Q#ӄH/� /kE��9��8)���:H�@}>.b�L1|�ͨ�o趰���U׮�*ƽ��y�ѴU�#ln�%��L+ݳ�!�e�QK�;�p�alO�1�u������5T�
��~�Ώ�i�(:�cz�ڪ�u$RH�$������
j��Bs=q!ho�(��$��x��ܴ�-�����J�jL��&y/�`���VKZ��6E0�K�7�1��'�XN�ݦ7�A}�p�(p��!D�sذ
�!�+?���͓2[��s��.d� 'HѲ�G5�9�c��7JqI��O���@�'�+��y���c�b	�z�%Gܱq�e� ���@OfN%��=5~�i�z�j�vR�Qƣ�J��n&>7ئ�����n�A�t�^U$	�Ҝ�%�콑d��P��y{9�_p����L����U8����x�=y�ڥi�?m1H��HK
4�I��t6Ckb? +٩�[%��F妏� �ܭV<ܫ�]��X>ˋ=+ݽwB��(�_rJ��Z�tQ=.Fy޻��1�RS��FaC;��z���F�Y�x������wlE�c�0>�By�������2~08���&3�i0�/�n�r�Q�b�dP-W��F���(w�H�JZ���hz?DB5�qyQ�)җk�/9�X��4�,�=��ls�5Z`Ƶ_� ���r->�>�X�-��i�;�T�nϸ
��-�sl?ϓ�*r��L��=T-����ѯ��b08�Ш�j�j����9�l��)�^�F����)e�@��g�[l)��s&[ذy>;�rlO��o`�fNW�X�K�qMd�IE���i��|���0� �'�����,�	�ͽ�t)o{_��y�H��+-P�+�������&	PAy8���j��:!?����>M�Q��L�����>�<��y��x�VA���R�[��B����z;��!�-�:���Y��W[��̀�_�z
���<����W��檰<����}��f�[M_I���}��ĺ2Dlzq\���kfl{����,�Z�X��\�#�8��F\e��r�Nʏ7����d1`�&4T�^F-��8a-^=�i�JeI���~��W�09T=CH8�l��Hrj�[� �^�,���찵�Gl�b��>L���ͳ-� �<P��ɑ��ju�M:��,�+k��Cm����"D>�@S�	�^c��Oq|�34����)j��:8PP�T�Eŷ�V�P�NH������x����4u���[ƶ�N֍xM��P��2�{���
�y��z)�L ��C�	w�y�	,?��*����3o�*�%C�{�po���{��.��j�Ͷ@%����t��o�`M��7�����]�)Ď���+�����2VY�;jR��Ԏ\�g
P�����5�Ь��;��+�pdF�I_�F������k�
�a���I�_ĵ��J�