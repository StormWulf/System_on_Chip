XlxV64EB    fa00    2e10��v�\��0X8��T�k��3���l쳅' U47�Wݖ,2�t��P��r��� ܥ-=�L|�6pa�e��bӠ&���qϾ��h`)w�aČ���E��jMk�p��_w/����s}���[M�A������>�l��g+`��}��'�������{�vl�r��9_ضfcM�[C��W� �H]��BS��e"�.Z�^�p��x����r�K��ۗ�H���o�w�z`	�:�]Qn#�n�_�ο��T$�%���Нݲ{��@�+聪����Os�n�f'�T˜�2�~���87�Y���Ny-ڻm����?S
�||ݻ=�l��H�ŵ߇�}�/(���@,�wʟ�q>M�w�7��X�h�t��<H�+�U!>�/QǮgeQ�
� ���>�@{0��^�����j�F�ÚJ���<��z�:��Z_�z_sꊥ�+�u_�wU��i6 ߤ���s%�/OL]�K��f�O
�݄^I7����3y���9}��wzqf���^����ٜ�i�6�dX���5�;����b���c��0�<Pf�Ǟ��<8�hB@��|�yJ��[*�LP����[o�o���~.2q�If�$��u�%��P���奔P������ޟ}+��ȱ^���_�Ⱥ�������޳��Io8|��5�� ���f9�n�/T�G��`�;�-��W�Rq�;_cۡ[�I�(�OF�li!V����l$���A���ٌdݕ���_1�=-�&X�� �J�0��hRAƆ���5�]������x���[���qj���Z\<_�=� ����Ynd&(���^A�ܟ��7�S׈oiN��BP٠K����v�?r�����������T������^5�6<ݕ5��y�y[�hv�L`�|�|X\Uv"	��A�̓�G�O��8���ڜ�����ā�I*SL�%Bo)x�-����%Q#�U%�~u�$��dɕ$�4y�=k����}�(�$�e��yy���S���n�F�|`RW��b�"�'v�Z������*_�ۚ�s�|� ֆ�fr��Y~��39�����S���8�f��/��j/0�S|TQ�e�����-4 zY'n��Ia,CC���axm|������S�36�o���)rl���Wp��d#1=�`�2w���,��س�,�f(U��.��d��-����S�]R��3F%V�qCݝf6���[�
��"81�:�D#`2&�vL۹QKv����"��M9hm��Q�+~���)��Y��0}��u)�y�"n8�ow]_��'��+�W�\X���+����Di����xX�B5�a�N�20J��LU����o+| 6�Ǵ%���4-��O_D��i�Jb~cW�D�)����Y65aH�$z`<��8lG@(�N���o����X��>jd	S�-~��Bz鶌!9��0�a��ew[����P� Z�|"%q�q�$���[1����V7	1�N�}[֌��+�83�&��:��fePņ�!�@>�B_T<��QS��Lb����5�v�O��h����WdT3T�yF
���?�yc���4�n\T��BSU(v��)�_M�O��M�d�u*�W@x��/q+�/��:Z��ٷ�PpE��0�2�h���^Q��N�	��a^��|��13�ǜ��߷�Z�=�8ѥ�&��9�]H%���	�D���ߡ<�R���	��i/��Wx�R���Mn��%�ud"Ψ<�K�2��J��<RA�*$+0��L�4�Q!����yY�$3���-�>�XF-�	��v
��	c��ɩ�t0������a��-�DQ̉K��z!�PPW����4��_ho���ya!�{��h~_�ݷ�E�;h=��b��D�>��o���$�~/{�˾=�e`a�2�4�(���H���\�s����n�s�^��k�o��Y�/6ǝMQ�L��R"�@�'�-�Z�Շ>�I������� x#�K��CB���l��� �cU��Ǫӫ�=��_�ǆ�{0]�X�y�Oa���l��@z {��`�n���iɷ��"<�zڹ\ǐD~�WֳwU�{�V��dӋ� ,��v\e2����π�M�H��]c���e;��:٪ݘ����%o��vlS�KT*���3&8�)OW��n��ئ/�L�s��G�D����"`.H�/��Z��J��4d���ey�IN�ȣ���� d$�m���/~ݼ+ Q??�ވ�0�U\��gT���8\a$V��ZW�{�:����*���Mp�����*��]��M�z����C�%����%P�x)�I�&�I���{�x �<�S��^�~m?Q<�ڈ��K+�&+��kպ'�����hվ�ea�0��S��P<�k�E��7��9�l>�K��?/���m����U��g��G�@~Ty����G��,ȩ)x�>��z�}W�p+	i�F���3'Qh����(���YpBG_/��Vv}́�9I��į�s[�A(7�3_��HYO�ٸ�v'�]�ώL�^C��w�d��雥Qt?mP�@��D�9+�����	Gz؊��$_A��AQ���.G���T^W�1��s�M��t"��R�P{l�\AC����DR�H'vUjZ�h�|KX�KA"�zAE�\��E��H
̡���׭�����u�^�귂�=SX��$����K�Jh*�Vi9������/�T:�Bk�Y����4����{�"��8�H���H�64��k�d)��oJ���]'�� �`��,G�--CJ�"{�J�s����pQ�
�7Fgq���ۊ8��P��8��Bt�6���lg{�ck����M<������W5����s�Z��l����,����#�F�f�̵F�>q��v��6�k�kU��1.���lHdӗ�q�=���Y���24^I���+���Ỽ�e���6���]P�Uy|��E��Oښ����$�kXr�>�wFFu[�o�o��;,֤���~QVp��ÅA��|w���Z�U�ݦ����������+Ae�`��5X���&�4��g��4��8�:����+$�!2�nb-j��zr���3>�?�j*
���I(��9� ���I(�cYbiMۍ̬=1 ���w�gm��>+�à6e��*��������w;vM��HCnT@�A/h��6O;&p��=����O���f��ڥZ�����&��o	�s[h�?g$+��5کQ+T�Y���l�P	O_*t8s�(������I\Ԝ!c�XR9*��q�}T�6��-�
=�9��88HsCU����l9�ë=	uɊ����w:z`|q�n��L�y��k"���H�j�	#J���v������Bw��c���ۣ�Ń��˙j���ED ��ۯ���ǚ5�|X���њ�Z� "���5�f�,M	,�9�}d��J�%�a����@6A0�}K�7rbtqOɊ!������=���71*�Y�<�����]��mB�T����	���$̆���b�)�-<�ղ����6͌"��� ��$� y;5Ə�tb!�64Y��~%�i{���b�����M渊�p�b��fV����y�%V!����J����^<��=���=p���u�>9��m�t-��d� p#M��Y�����S� }��/�ľ�o����E�1������n"�E���6}!���$ڶ)��j��2V�:�vO�O2�_��2.���ј�vN�Z	����/�c7ː¸,T���5Aޙ��DO��uD b�(�f3�?�2� z�
��"�c�U0k��1�J��]�����Zq|�D�+8��@-8��z�|�V�VE�m��ތi*[5~��ZK��M3�o�9�����6F
3�{Y[|�[�`x��ب.
�WK�� ��Тl?�>�!���ѝD��δ�{Zj'u����	r��zA��ބޱ���H�̘�������c]�~=���)J�[sk�+�`UZ�]E�V<Qj��Sd��p�G_O�X1�q�:�u�VY��x��˴1O�)ɲ�x�	4|��S��]�0]������Op����6�ˍ+͌����w���ÁBu�F]&Y/�Í�<�0��0+K�⤍�����-Yn����&»[)!~կUP%?q�'5ȵ�m!!
�f<ҩfY��M��yQ��w
�/����uѶQ���e��iM3ܞ�Fy��+u%Ͻ'�>;*���l���9�<�5�\ ��7����[�è��`#����🄀\2�3ۈ������9�ê�'�&�n3�,����������c-t�(;ȁ���d8�+:�g�e4ݎ���GЋG�ҨȃY���&����7�p��vI�w�ʆ�Q��[(0��13��z�FT�q�V�K�`'�J��2����a��:`��f1x���N@�JƐ�- ���dZ$v����� V��J�b\���+H�CH��s���t�EA�&X&Q�#&�n͹���%A�G1�sڜ�1�t60�m21Q�
�/�����MW�ɾHJֹІq�<U�@R��)|ôM3���ż���@���W`v�BE�\����o�c�I�]��6 mxHU�숏�^g�,��!�΄��Ѽ� Ӝ �E'>@��
}p �b	AM���'B�X��UC�+���c���Y{�֘d>U�4sE�O�)������}F��;��K}�ګo�)���Eԡ�Җd�����4�\�u��)����`T��+|9R�z'���e<��]���.N����/�($�E�Ho6�y�?�#�-?����8���)\���[*�%s'�;s<�?�p��QN����ͫ^��v�C���]L�7ULB���P(��[ �l�����o�oL����Q�a���ܛ�$f�̽2�N��#N:)h��.��-^O$�sDQ/��C	D����}0��y�N��O�=e�B���1��cFҫ�;����F+�����|Ʈ�l5���>]՗m|h�l��%��:����`ag��z��c�@��yN.O}'9�ީ0���WrOɧ�7�	U�Q`|�B&,�t�[��:s���$5�����K�H�
�>�e�W��aR��Re��W4�l�<�T`��6�5���9c������2�0)�G���5Z[�3�24t�/��e��3+rH�}oNM1An��[fe�;�-��&h��zw�1`\��k���F��ߝc�P���W~_�����>J����S�I� m�ӅY���W��|
K������V_��on���"�E�E��̨�MB�ѯ5������;z�;�ٞ�[���X�+��_��kn��#e�POWk!��;Fȳ�s�I��/e[�?������M�k�����GWO])�g�oQ!L֛�lq�/�MIB���ɍ� ��j$w�3���Ѡ�0���q���j�g�X]L�nn���3"^��!D�������P��ô�l)S�R��^����t��HpnE�=!�.��;����O�	�-������8^'V�"�y.�Ӌp�`����6��Ql>�>o�����P�.��u�����~��{�>��3#t���J�%�#N?��eMI,�<4)�_�r�~&�c�����O� P�O�ԯ�/��'�_�H�Y���{;i�W���((e�_~	��e('!�
&�bտ��e1�L%ɉQmB��+���>7�C	d�9���q%»��E�92��U���3V��/�23��@9��O���H�H��L�B����3/�f�E�Y��A�{�_�����^ڊS�St����X�N�׃`�`Ev��}���>��`q<^��{�{�nT%{�j<]N�O�@X�<�s���bV��V(|��dw�q��1�E�3'�+�u�="Эnd~���ua&��L��O�Z���b7���m�� ���k�����>iiP��`�i���܅�#�kCV�/�g�[x<��E�����F�W��mA}p��X�
FL2���S�(�l%#\&�՘�'9p*J��5��-�i�����TF�$�eωt{~�gX������%��nܞ�T&A_z����`����WumT���8���أH��2�%1M%�8&�9p��P�YzF?�ƾ�S�����7����#�:7�Ɲ5TXQ���K���YLw	�S�*���tb�P���`itg�e?�-��<F3��mqa4��0�$v���+�r�>S0Q9�j� F�����U0�Pj㈯4��������/��T�u޺���,$1���=�R� r��t%���k�÷�e�B�����4|��r��G�0���hjP�ơd�W��#��X��=������	F�,qU��1�B�d)JcюkA�n�k��L��\|,�)��I ����J��N�o���O ]u�zy:��_j���I�
r	w�-u�D��m��MG&{�<dKޝ(�B�F݊?6z\�2L�W�z+�同�zS�A�Jh�f����3x��,,�wԱ���CD
�"���fQm�}ls#G����xm���~�6O2�K":d|M�#rBs!�{u|�9���D�8���3PKۘ��B�,|��)xw�R�L�a��~��F1���o�Х"=�>�zqGE��c������k��ϱ�,{"���?nP�'��Ʈrd֋zR!-��7~�D=&�Uu<��8r�3��Q�}ހ?f&)�����b!^���� �K��+��-�v�C�D�*�C�0&���H�&)�z�`�I�R�[��ؚ�2	%g ������ǤΎ����ۑu�yq 4�����ۆ�Z��k�M�����&���g[1&�ɣ��N^=�h;Fԫ~G�X� Qj�`�9W�R0�C�{w�bOE5~�ܴ��DQ�*�)T��R�/�D���S(�c8krAS?��$$Kp�����Tp*�ʹ�@�a#R�\�6a�C�d�(<x�
g���FX�����Z�����SrДyeU���l+xx�:�S�̐��2QJ�ᯰmc�(1ٯ+�Y5ǘӸ}�oΕ�Cل�_$�E� �!#-�t6�3>w�I@I���ŬM�*7��1��o�J�=&X�Xy��̍�lo�WBf���������]�-G���p��7�v��-���b�ϙ,?�b���EJ*n�>r VQ�a�ֲ.����!>IG�n׮VwtB�7+$;C`���@��h7	^�6�A)�d�e����a�S_�	+�k����vh�
s|o�Q�L�ux��iы�[��m�I�Z4.Չ��]�I��)j6.�E�O��g:Ky( .�ȋ(����,�f9�r/ ��0�ۢ��L�@Y��EdL���{�7�V VH��X?\���2
���z��J�]}q��J<�,�\�ǀ�W�3�[�|i7n�FF��U�1������+��K���.'C�����ڹZ��Q�۬;m�,V�������j��V�`�Q�I�Ebmip��$�.l?Z���r�|�<ˎA�L�����7�c΅���@�yl�d����Uj�"� ��FٖV��2�i.Zl&܌<��h\��Z:c�7\��-e(�v��3-Pʾ#T�
8�S��^#�-�� }���.p�<#:�-����(*�w�@
K�m>�!�����@���;�+�t��GaZ"�&"��s��g#�Dug�샀�tA$P���ʱ�37z�c����:O�j�E��{f�g���j�� ϟ�&�
���d�x 2`p*h��F�0T�_7�
�>��v#���^���ae��d�A����?��n��f�}ˏ�S/������YZ_����(ޚ 
Y��<j�#"�~͹$P��Ƥ���,��/ ��`��8/��5m1��}���%��c�}�v�7�.�q^�3���50�f$��R�-�7#��Q��<����2U��	Z^�T��X�"f�gN}_.��2���;��qԕ��N�|�����J��X�#��Ѽf����u9��(����>��3�v/�زE�[��S[����f�w�3�*����2\�yOSCD��FH�.��l�#

��[���r; 4��h^��Fܲ6dW<&���*e!��k�b'����Q"A�~�]���/���ҿ�r��������4���� �;�7&Dg�.&�X(c��\/� ���h��I���:~Fů��o�5w���z�E���'\�<���oa[���}y�yvp���2��2
�Z�:��*"�T�\�D�p��m��>�]^��à�{@<ݩ�T��+�,|��Pf&��!�������X�r���-�<��7ϡ�sYt#��q��o��nz�z��y]��g�����
A
�����:4�F�U m��������ٯ]6
;W�I���,\ϔ��4��A�+dX�c�O���҄j���vg�������ñ�B����d�k��9�q2mt���0M��^j-ѱ� �=g�C�f�s��q�,��TUu�(��^%�"�#�|��b�֖8,[�&��(�+�·ɁM��������FFCP��=2���]����E������9�
B�32(����'�����y�{����xt:�@�c3U%0���J%&`�t�4�sKj!h}���}%Pjq'�#t��N��������K�g���,yTt��u�cpT��w���hN��E�#�G�XI������!���]7�
n�9�'��u����Ľ{�3���G
?y��|]<�Z�d�~J����n�h@�\�bWM7��'���)+_����'�V;���'�e�	�fS�Ժ|�%E��X <�`BDb�Ԩe�=�c/6]G�B*��F�U�a*�-�8@i �Vt}�����y#�]����-:��sxSof��lGW�ٟG3C�:��X�R$�.]˹�!Ycʮ���L'[�'Sn^�l(�M�fD5������d�k�s�TT÷�l�u�o��ԅ�#rA�G-�����FAw�������������y�sڝ��'!���K��|&b�1t�	��/#�\7Ҿ?韗��
��6~h�&~!�.�#�5�
�b�0�+�bO��v,��d�Hڝй���?$��M����H9�}5�(Br�GZ��M"=��nԤ�0X�~��#`�[�!�I���=����~�S��	��vU�F�8S��U_���΅vԥ��=>��)v+t�e��e2��"��N�o��v�����5��a��#RGY������,�ԩ������T*�����@r]�m/f�+����7��7�vm����� �!���D����c�E[�w$^h���igQ��Ξ ԭ�2\���^W��#`�grl����L4�0\��(v��:�����M��� ʪlA4DHc:a�ZA�'��	�?�g���1�Z�œX\�dI�����DО‚;�Ҙ�X��m܍-;��˄�:S�,�w��ps���"����C��M�'IǰQ����ڧ-�g�߱;�p;'ˍB�U޼��kP���	�KHX,"������jXl��G	�I.s����T�_�(�c���ӗGwv����=���3B�����M�Fɛ�?��ւ�:Դ��ގ(mN�����=.� �p=)h��yi�K���H��Y�}-���ȩ��YĳV����
�'F����G�Ibe[�5�)�z�Q����!��Gg��=L���Q�}��<[��7B��rAa�=��Y.KAF���-х+��(�EL�e��H٬?
��
�t�^��<ӷk�o�S�e�Z�|�qQ�T�*P���,�^�����7&�ʅ!o���^
���0��Qj�ҥ��ZW��ݿ�NM�W����Dw�R�À'�@	m7ĲL5o$b���$5k57�Q��,łef#�UIМh<��=�z��!����2K�̬����
cܠ�>k�,�Y�7�@/��` ��.H�֒�eA�(�i�� ������G|*������D�L�,�܂�p����A!��;[���eK���<<k���lf��2	�� |r��	8��l�����cM���T�]#�N5ʍ�6�M�����\d仦7�n���U�������3D9������������N�|�Ր>��8+������i�� �ܘ�];KT�M��}N@�+�j�Y��������=�1�_�`�`��[����H�扞D��c/m�A�)ls|Y(w�8cdu�gѾM̖U�H�d�/:����B���D�B�h�ja�m퍱�;c㯂p�C`%��>�b)��L%-��b]L���~a��1^ベf�:l�Y�=9����c��. ZUO ކ|�%b�-JJ��L�}���R3�s z,ޛ�~xt䨫�D��@��W�:�ץ�/�զ�][�iV�~>�s�i�X1�2P�J6F�B<��pV���`�IkQ���S�8�yf�m$��� ��\ĭOڟ��{�����O@S��܏�nr��n}q�#bR�Q0����@[&	ؘ�~2/��ȷǥ�*+�;�y�W���g&Qy2�［�(����l4
�}��rrP$/u��W?�j��X�i���~0�҅t��Lsz��0|���A�/����^�;D��Q}�Nm�n��vU�����XO��yJc�>�s��v��oc�P��vh�0��*��g�)y�gM;S�߃�������B�w#���(�!Q����g�����wg�ed|I�(۶�L`���	���lyR��B��w"��*XG��>d�C�g�uE��+6�nN�V�LT��:�3���;��Jcq������xe�WDn���5}�Z��F�"�����1(6|n
�CPh`�D��wUc0�3ᶈ�I�k�n'�&���$SB�<�\'a-`��c�q��Vj2�����9�zZ[��͙i�ҿ�/�x
�CQ���_]�M�+��o���EG.��%'�F��#��Lg�%(a�{e+���i.������m�j�I>p��GXt�	1���w�U�=��u�3q��៼s�_�蜑��E����HX�Y|;����������<��:����#��bVQM"�z�(������ww}�[�Wl�B�l�%Ȋ}� �/*��ʱ܊���%�A#K��F�e�`�aek�K/�Z&=/y�1�U���a2u��8��V�-D����(�e��L-/.'�W��s�=z*�6��\���>^���b��\�k��}��	KE�;$6�6�q/M����4VEj`(��I��el �<]��r8��2m#�#�*Z�	�$/��^3#4�l��A��!���#��#� QK۸�QI��^6U��3�a<����8� �N�=Z����ӺN���d�U��q���@U�	�_��C��\�f1�t[Q�.���Hc�uYP@�S#��Nm���-g�BJ�8
��=���КW˝�ײ�W�1�{�ڼ��;.P�H��Q����&+*�����_v�4[��:Hv�TpA��_C�	Ks:z�W4YP������p��3dvxl��,�$�Ī$Ð��:hnm_̳b����r�d��_y.����9���X�f���Ң�HeE>��[v���u���:(g[O�-��L�]:|���� �хq���`:��� ���&/XlxV64EB    3f4f     b30)?�,B�΄q%��̻�&�_����'���e�W������ɝ3�F�A�=�t�oӹT(E.[�R�<-BD
Q%�&�c��5�{*P��Mn�k�f+�����ݭ�F�p��IM,���n��	����i
��Sa/o����Hصs�L.4������&��)�g��!qgQ����J�5��aj��W�aq��� V|�b=���B#�G$-ցb�T�� ����GMgc���-�Q�E�Z����U���:����^��.����ֶI(+�6^'lT-2i�g�ب]eL�J=��-��Se&݄����*M/dD�[��G�R��a"���������q�o�Xހ�˭��m#�K$��y*���Ẇ�V�R�S��/#h��@�C&	BBF�t�|��@P��@�[Lj��t�IR���>�my�l�)$!���5�.�_�:��\;G�B��K�y��Wɻ-����J���w���ۻ�[�{��OlU�xr����<��mI�||�?"���������nx�da��E��FG[���hL��{�t�IŪY�t�	�.g�/toqZV�{.>|�,��$��a��#��4��}6��-(�{	
� ��5�Ʊ*��������$�W&��:�<�e<C3�O�?p]���e��s�e=icu
E�nΦ��5����BkY1M<Q��(�5��*�BǢ�r[��[�7X0�(פ|q�,���9;�ԊC�� ���d�LZ���F������`�����8*��f;0F act�����P�Ns� #�_2c϶�����$W7忀4]<!z���i���$tz*�A��
�<5�%7`$I����:�Bq�W�n?i�o�Cv} ږ�ΐ*��
k�qn�7 �,�5���4x�h&-�9�D���7�L�4�4�
ꄑ-��}��	Z��q_Pғ`B��g�5��m��/�ȷ8�=C��:�8�}�;��g���Xb��������@��=Y:��z�ΥP�O�������3�n�"���z↸tTt3c�&פ���s��i��(��֞ �[М�0�s�8E�sW(�����dq;�hso���Kf��愫����$3)�㈺(K�a�۾��N��̑5%K��@N��]�E�<��]��QK��ԉ�T�Q�NU�d4����:���e�{�H	c�2J���Cc�lװ��,���oR�ѣ���4}0l��Z"�ɩ%��8�Ժl=�e*��B�+�#�*�0���RE�����*�\�Y�gE��
���w8Ϙϥ��D��JCn��C��B����#��<�_sT��p�����xW��P�$��d 䕓_~�9+��]
����b�ܛ�Q���L#�*xr�caܨ�m����B����~���� ��G��!�8�uig2J|�'*���w��<�}y����8�PԤ�ּ\i���M>���]V��N�F���6�s���)6�+�i�ٿ���\A�8y�=��Ҹ l�,G���A~��蔑~���0*��PM���N��yu�ؘA��~3>�s~�S�ɟ�V$i,�ahZ�X����aΏ# !4�ZMh�塁U�e|�w��5���R&�@q<�i��Vx('�-(gSp���8�k��-�2Z�ƛ)Q��X�g��*'Qj����U��T&���̀�H���mc����;��@�+PS��\ y��������;>�}2�J��p�&�0�F�N+�b��G���k��:��18lb�8[,����[�A�s̙���P����'��Φ��@�`��0�ԏ�f�4�Uo=e'T����ߒ>6m)e��l~&��hӖ�JQ�č뀈uDBX����O�bF7��A���>K�����]�h��qt��X�Dg)A�*�۳bQ��:�H�D�>d�$W��E$wE�θ�𦴤G�6�H��.Ӂ������N��3�����Ȏ_�F�l��9!��2�&�,+/����,+�'L���T魐ɍ5t��n�U��t���}�A�S�"祝s�-��)b�k rϕa.O.x����XMRD ������8V&;�P����ӰS}��{K��0��uVeH6�蕾�M��
Ł���@{����ة���p~<no���q�X��7f�5��8e�L�nY�b+�V�!oݩZ��L�E'ǔ:�gIGaՍ� �<��X���\h�`-m'c���^}�y��_)r�������Iz��*[�B7f��Q�R�V#��0�M�ʅ
�^���P�@�zcɹFM|x�I,�6��a���J: t/]���^@���:D]��E�pM����Փ�Ö�����'	X��n�u�
���7����Rȥ�T���ц��D�KCA�ꔃ�6$��&��g;��N7���=V����Wv�d~y<���4�ߵK؟S�8	z�=�+j��k��E!�p�X�`Y��;������u�=���V�]}�o���ː߃�F�;��~82�H�e�r��χξl=؂[��ߦ����&���4;��9� ���Kx�_����3VsRWC��4=�	��>@����t�c��;1�AY�YL�ws�^3DL�.4�(�I/��ͣ�Qb�-��L,�`N�Gy>�>bu�zn�i�b�#~�*?HA� aH�����4`zl	�Ⰻ�J�ZX��B��m@�,�}�*��|��3�/HNm֐��C���sG�V0'tE���Ybj�6!��)5�����#��Iޥ�.�m�����)n�,�����U!�~�n^'N�c
��u��_��~<T���#ĭ�E��ӿ��