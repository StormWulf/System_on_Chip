XlxV64EB    2b47     c40<ĘJ~�3��=�D��`o !x_՚K�PL[��dA7�0�`�=.��WS/o��T��\f��Q�+9�ػ�TM8��2&�W���lsL�A7��WZO._ �2����b�l��R��Q��T�5ӉH	 R�4йOb��u�&�{hѽ<��^�-�c����?8ʷs5�k��`.3�>��UюU��g��ۍ+�[�Vv�+��f�v8�/�N;(?�����	�ܕo�į���t�g��v��NzW��U_��y�&ƈ��U&(���,p賷<��3l�����Q
Y��Ons��Ꙇ/��gj��Z/�3�ő��Ө�]4��J%��\��+ӡ��|����xL��'��� �"��y}��	�%4I(����~k�6Xܒ������Z}}A�垓Ȁ�����ɪ��P��� U�
�������a2���Y����UBK�Q:��}1�Pr1D�y 8����<�e�Z׏o,Rjmw�)��B��ZY=��:�����,&2@h�ܫUo���~Ce�_����0��N�Z(UC��cA�+�E��At�NwZY�Y�H.���vY]TCt���a�m?��}�D�2�+�2HC��:����՟�.�5���.޺l�  #��5=��/L�:нnN�!I}�1�|�H��f�h��w�t������q����)pf߶l��xLXm��u��E������Bk�L�{9o^�)���w�[����uuﺭy(|�%D���&8�<Z�t�r�Y�7pf?֜���������i������-SN�`�f������b����j`^w_�N�����ek��d,���`�����%L�)�*��R+�='��h��Xء>�[D��O
���;r��1�R�?��� `u 0/į?[��k�ي�� ,^[��L��,�+	��Jk�՟�oY�b� �q\T���gx;���!a$Ebk3��)^BQ��F�[�"���į	e����0%� �N �X�!ԩ�I���)��0�TG���c3k�K�)�~��>�/��p������38
Edп3t�eb<Ö&�J��J�n/�m��Y��`0��.s��;�aJ-H��%*D���A�(1�>R=0��a��^	J�Ơ��NSw ��@Bu7Zm����*�r2-b�K	��i�U�Bl>�qHi�$��Q��%�Սh�
4j�81L�����;�p�́�m��\�sJ�Ng��~�`+�_vc��yĉIy05:��tr� "v��� ���NI��5��ZR:�gR/F2`$w��� =:���m�dL��f��n}�↥���7�uAC�;X>T0y��J��;�w0d&�v) �ċ(�yCjg�Bm�r�OFU�R6�1������-��lE8�u� ���f�;+��N�5���۶�)פQV��e��bj�iQ�[b��"����lJ�!���t�����xࠁ7�a��=�/xKf�ɖ?�.9)=����Mh�8�[S^Y>l���J�y,%���>|`QP5���Z�'JH���ƴP��ū��/v�&��<���/�ۺܘ-�/��N~d:oV@�h�H����d�#-��/^���u��L�q����E��� k;�� ?��XOAp>�)�w=��Ҏ��0���"F�~It��[�������`t:gi@]tD������3��mҲ�Z�S���C�-�Q
��g���o��#)�r�?a[�L�r�W�t�F��L��ep?���R�QR�%�I��@x�H:��!ݲ�UQ��<��dH�ֹ��7�������q���U1*�B�p!rA�@��D��M�V�6;E|x��*)9^\sͤe6�� �������O�S�j�<�������"�d���ڔ:Q>fޚL'���@�Ȇ��֜8���뛗S��L~B�V�zUMЉ���jD�Sc�E�?F碣�4j��A��;(G�ӳ��p�y��:1�j٬���E%J�"��6�P�گ
��v��bR�ˬ98o~��-2��JE��!�!c�'���]���шokۿb��Ii�!��\͞i$�?�h�|g�e�a��@w'7n;ˁ�����E����H�����9�/�s�d]��&��,e}�H@��=�\�� ��<i��&�V��U�At�-�74�Z����k8�����b��'��-/m�Ql�3�s ���Y�ތh����U�I@�;p	�ߥx8��A��\%���~�r`����3�Z9� �V��2z~��d�Xj.��/� �9.������v|����!���E��jRN�r�5q��xR�����B�����8x� w�'t���W�gZ�q=���2�!���FU���
��S���!ʃ@-zv���-�`D�1���c�h+����s �p_�F�YB��%��܆b7[���Z��YƁ���{ �D�Փ���m��"L7�%yIP����Q�O>Z�T��|\�s��!(�?:^5(��yY�ڊ��¶�DR�����Y��ўᬥ_+����{\t�O��vgo���6��?{z��:O�v��퉥��|���-=��7|�� j8nh����h0%S��=i4u���/f�"�CzcE ����e��I3���^��R�E�H=�97��w�>����CW�p#J�� �6�r�Oj�q*wk�3�s)�x��L���8_��:��(\>9& ��8��/�Y�V!�'v�O��ϟ&���O�KWv��~����*�gT���{�k���l��yCs'|��a��2��u�NS) �Xa|��J9��=��aL�#C���N@�s�_'����������'L�U������o�GX+Qe�ֶQ�z��XÄ)f
}<�m�J�f����1�=߃ȫ@��X�R��6I�x�A��$��vO  i�X�k�����p7�%�Ƿ<�+twg�j��ӾL�]vb.��/�ew����5�J���}��1�"��FkJ��z�jfE�!�a����;�[Oн�RϘ��[���= [���t��vv̲���b�Hpts��S$r]��%��<]^^y���c
Q�Ր�D�-�}-�XL�;[[�f��p�!�i/�}��d�ٌj�H���;%!:�