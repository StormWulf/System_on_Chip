XlxV64EB    fa00    2ed0�#��Ҩ�Rյ7��;�̉Y�����d��Jc��q͕�����z�`���{G�!K'����Mh�����.��R[6
��k�2y�_���[�ax��zY[i�rLk�<���S�d�	�ҳ�q�V��G�6��%g[H�|x���u��]��/��J�r��:,TR��Z�ɗd���>6�A�|��m[/�=�7�Iٝ��O�sʙuA���iN���4_z�wj :v.����LJ=�(�䧒^־��J�˝�y�/>�D�I�p4�e	��C�C�S���ʚ*����W.e���R����58��0�������>���]��I�f-t�l��Z S�����QM���	�i�Zӕ�4C.TM�_y!q������"<�{L�^�_ }䍫�/ԯ7i��S�� ?ˀJˉ9�g�ſ�;Ҩ �i�������su��1Y����(`����g|P��VL9O2���T�v6� ?�\t��1������O�~k~0L;�
�[o	�8�K����}Ix�~%8Im�?P�T����>ē��6-"�O��:ᅼ�?�%	�{i�b��x*�J^"�|K0�wđۀ���3F@��q�����*���͉yf*+���`�6 �i�Q����,���Y��2MS���Oa�{���Q����9���ޛx��n�"��k�1t7�ɪ�D�Y~�������S&!'�d&��;��%��D+5
���U��a�"§�m�	�<���aT�%+��lv�y�1�P��Ix���V݇#����N�t�r�(<k���@X�}[֧~�D�Dk�\�b�M�w<�������n�o�*r��W��u(j,����>�lٹ ^�D�I�Q&n�Q1�IOb���k�m�n	rV���=�wO��ul
]D�;�̄����P�@2����/yo�Ǜ9�	Khw���HC�HU�hed|3=~*&b��|<yy[E�����f���1#�
��"m���0�i��Hw��u5*;���cMAtA$�)��@]�� rfTk���Cu
��P� ~Ѷ����%�<n�,�р�8��M}[d��恵�[�+�uI|��H �|܆B���(h|�e���L��W!	�a3�n��q��o��V�:ߧ�{M��36p�M�n`�{5����q'vvO8S���EB��c��F�F�RڶqџlvP�*΃�カ�j�ݔ&l���v��Jdr=�G��/i��>�	�v�-�5�����	<��
���J�=dLQly����TFSal&�`���j�ŷ��G��E�B:�O�t*��G� DO�UUF|A�!@�n	���/�Q���o������ߜճM�;�Dr�� �"�WҸ�b�9`|��Ð��Qn�h�26QlVʠm�����<�!�Li�o��oc�+ޖ���5۫S��<�W�%����"����q!��Oh��^��� 1m��*�!�=�̓6q���>��ž���;.!���A���&VQ)%��ɲ�X�u �S1��n'����o��צ���=����Ʋ��5*T�7�.���<���8���Ў3��5V.X'�W��M ӑ��N�Տ�"J.E��.p�u�̠�W%��>z�Y{�sԧ�	� S�b/|r�h�uf�Hv!�^r�s�FonRƄ��w�p7����{����8$�I�}r �N��+� A ���?U;hЙ�m��4�����
A��d�j}�PU�i<��A[�iMB�\�@��kP��}E�\�l�Pb��w
ʀ�P�{'t�0�:�;�.��o�O�X��	����rx�Y̋rR����ٙ
M,2����a��H5QX{Y�J�"�~9'����Ҷk�ca��F�-/r���oS��~�	M�Xx����\b�ޕ2=����������_�����y=n�;`�G���pVrV��_̂?cĘ`��~Hd�ڮ:�h����p#n�$_g�L���[����%��ńX��������k�+A��l�����,�B�L�L ֩��*\M�2��R��U;<@q��xJ�ZhG�CGa�V��Y�hmzu��?����-���(���?��7��VD�#-m@�.2q6���(H�����c]d.MB�nF��܋�����)-d��E�7	rxm�da�wJ<���Ԇ/n�����9�t��� *Wd6����Qp0 �Rv�x�/T��?8[TwqV�3T	Fk��'R�%��t����/�Q�����?X� _��R�@�0�\�
J�L�]���������a��v�ꨄ��^��G��#c%���5Y��nwb�\���
s|������gC]�Ey�rY+�|q���:�3<�+CX9�B�+4m�9��)�#q\/�zi�m�)^M�g�c��)1<kT�VL}�c���8�'}��C�{�>�[E�
�b���i�gːx��n���f��r�.{���^vg�b��J�O��SE�C�T�P�o�Z/��g�[��ل*Pjle��D�ƆBx2l4��kx�3T�L2��G{��b��Xf4(����3�.�h���@��zK�/�G�"M�����RtJ�r�V �[Ӎ6Eu�����0]�9���G�tP&~馧�"[��n�^������PYj8�bX�8�)��IY@*�nڶ�N3��ɚ����$��[�;ǝ�%Tˁ�[�YA�4,5��b��YR�B�
�k����D�c��ù�p U���0�g��*�`���s�	����,-3���mǮs���#���" "����+���z�l����Rp�h�ߐl�Oв�Z?��ۗ�%�y���9�Hݮ;�a�Օ�{�(�k�(4�o~�oAv�4�,�oJ?/%����xXl C�Ԟ��HJ֘g1)O���H�H�(.�^��{h�Κ��,�f#���hz���"K�å~�HE��r��1-Id�vW���X���~��!��O��w���,���U��^�=6�?�2J �n^�W4s=�W-̉����d��,���
v��9h���񩷬a�-n�(b�rg���H-G7P�xĝ�3����/�D ���sf��^P�ye��Z���5�P��f7��W���\��7fT#B�Ւc�eP�WWje�K������"�����	���TV���btY��xط�EٗQب�'��Q8�W�@Z��G_lAD�P�ǉ*ɕ�ȧ�jJ���ya3���d��b�7k%�����
�3�Í�)5�q��Z��d[䳿�;V�1�/�.m[�%�R�y.�D�{¦l�#����T�(�����֍
D�h�#�sݣo�Dl��w�T��D��S
,Eo��l׻|���h����B�'9�o��vk4>FX��SE��K�V�qi��*~u]�jH̀��iHϐ?�>��Y���KzH�^�ȋ��IC|Uèdǡ�O�<P��TX� Z�.�f�l�m&���h A!Y��©���?
O�H&h��r�[`q�%,׵A�6u�����7V͊�]P��< �>��N�Շ��/�Yd��)��Dk���q*|?�m���L���2̘��2��J��@�du�����B��z�E�@�_�k�!�s�?��=�h�[$��� ��H�?[��]Gi�����a3����ײ�~����s��Z�Ie"
��ܱ�6t���~?W��*�`㱠(
�y�X�.f�������.�(���mˏ�ŶN(� ��^�͊Wq/C((�*��_�_�p�8,����<���"�̠�yq�j��H���m�
Sf���=�=x� ����m�3�dj(+�K��Um�B��K�T4ͅ��3�KLn��%�esx�W,xT��g��b�mm��W�y���YK�9����8gpE���R����q��Ř�դ�o_�"�NY돘"!Z�%&.Q!�������+��~�+�pW�ŢH����j��}f��vÉ�hb6-�L(�c���p�5�O\�;�3��l\������w[^%^E�1q15�\/�NNn$�<|�&���.o����(��R�Y.<���DH)^��M���\ն20�� j%2�.;y"A�j��$B�����=g�F�jX[Xa��+1�dXYl�|� tFB���[���#��Zp<�[�n�(�`�\]BqP������}^���.�)���PE)a���� ;P��L���"7,HC�;rKƁ!2�x��3�Y������p�
��
�����@ p�6�%��w@ ��#�`-J����WxZ�S#-[d�p��Wy�ol)���Y9	JL��W�D�&T�Ѩ ���`��VU���l���>`�Ğ���N�D�^V6�������Z�0ʥU��3�D&�n��lsH���ޢ�:���`Ҧ��]R����9�����%�Q�b����?���z2�bg����h�Yؑ�) D{�������*a����i������j��f�56�ޒ/��aD�3��1�E:F?�ŋc���;>��冕)��0k����u9VjK�:�+�=�y���2�\b�Q��wg�4''/��a�)3����ݭۧ���Rύ���,����q=?��%ne�<�?r�:2[Q��D/�C��e���?c�+C��N'���eS����ǔ|J�uh|�)hKO�k���"�N�:ȃFM�?��`�8-;�(�=���S����G��^���]Y��;RG��b���_bX؅
��)�q��g���9>>8�!�+���z5���y*�d���G�Y�p��m�k�-�Nc??7h��Jq�U���8�q*�Sfq��ݪ��=A"(k��	��bGYj�C*װͤ��NP�3��+�z׸��gV&���}ڝ�!.G�Ƹ���7��o�ds��9K�h��.�4�<�t��cV^��x
�Bn���G2��q6��r��'�0K>��b�������5�a���n�2T^�e-�i������-������������~�WZ����no0\9�0Y'�����Ru��絖�W�Syޏ���"�kw$��j���1aUjbeG�V�d*Qu�;!��f��N�TN��*�F
JB���;|�t�x뼖�C��c��c���^��{0�S��8�@���y��3X�)ߍ���Es���u��I4�?Jkq�=nF�#�z�,r�B.��g��Ǫvj���Xp����0�u�I��)L������7�QF/�"�ܗ�^N�߅��pA��x�R�����A����ʚ��u����AU���"|�Xe��p��.�T���z��y;�U�0�+�̾s ����V�*�o-O��l����.� ��ʤ{�����wTN �o�P�w���Y��R��X���^~q�%��%�
^8�/�K/�F"��Ҭp���?�	�0�{���r�
�g�nj_���M߱Z��f����f�Sh0�Nz��A]���O��D���v�
�Ե�������5�Y�}�3��&?�B���Y���z\=���e�`?�HI��-~	�+��s��� Τ��{�Ļ|�e�)R���e�EÛ��DA�HX%��:JP<�27G�ߚ-GlV��w��+��l��S�`�%D��s�Y�?�N�0����4�b|�q e����ը��ɘ���fB4����u��)7U�8�Ϛ$�����/��^����@Bx6���%��k�Ir�ɷe��q̼�N���S�Y��ةli������iD���p�	���o��u�6�X��xP����UV��+l��z}��8XEO��������]rȢ1����U#�51�i�ʴ�	���qr~[3P:E8���j�V��i]�IJ��9吷Z��T9�%�w�?��g���(�$2�o��UJ�H��{� 1>Z��_�z����*<�)�| h3�O�:��7��A!544g�9P|��̗b�a��R
U�l t�-��#^'��s(���c��U��:W��m_�r�O��p��C����kզv��q����xF�%��Ɗ�qt9#j��v|G'�R��S%��,���,L��� la�ǜ�����;K~}7��^i���V�f�%���<�
P|S.\7ȏrf�J��D�6!�,�=壏����I/8�x~�N��ꉣt�ܞ* � �$��(*E���#F H��[{[(�l6�X���cn�>B�&�&o"S�̝C�N�����{^X�X��Lt���5�Z�27K#m��ǘN� d��&b��!��!��E?�����ǯ��y�V�(��y���.���0�X�+��ƧFs�`�p*b�z�+	L�[��#�rT�{�_z�6K���w��h~��D��Ih��-3���4c?��e0���I�M��=�;��]:�>c��o�q�JzV0W�ؕ��q�f|�w�O@�k�`��B(B��w�hi$�s.����s������4X<h+��gG������_���W����Tl�bh��*x�r� Yv���&�1�Y�˧ʹ\0=������⢛`}�6>�h��=J�`��n�V5�*��n�>��pѩ	tm6G?ĦG�L�b�X0��?��Yp�d(���pc�$
=!��m@9_uKZ=��\��FoPd'}�YVC�Dd)���v��s�o�S��N��������Vy��-Q}��Wc#dQ.���?�;�J�+�#�F�=[����e�L0_�fk���K�z밤d���\C��y1��#h�́sGe���7�^Ͻ��DV�}Ǥe�/D@}��Q���Xz~$}gn��ʽ�f���%�L���4���Q�`]�{Qo�6D(+}+߳��g�}pM��\ayq);{�&�W���G�}N�@Y~���}��
/"�.�����7o��;���a@{���xc���*{�?�������7�R�:Pd��?<�+���9@mĊ�#M�jZ9��o��ut��Q����1�j�xD�ME���J�@�JK<� ����8y[�$uoW.כ����M���z�K�'[}6� GEpǠC��)��<�U*�@�Ŭ�����v�*�+%k�.P�o��A��3���H8����$��u׾�;ITQ���D�\�������1�05�Y�s�y��7��$Hu�m}[� a���j �6�r
�ɵ�Zf#�#=.�i].��;����f�?]-E�,j�nE�����Z��+ʱ_-��]RZdj�&���KK:9�^��xx�(~���2����#�B~le�����O������p�.������]�nq�W�k�u�6��{��U������I��e���gǢY�y�f�O�y_�D}�����
_�â�$���50�X�+�NT���+�N���]0M�~���$6=���#Ŭ@i���5���@����t��Y	^ZÊzf/�,7c����yL&ap�Xfʂԭ�7��Ly(�f�k5���!��+�Ɋ�z��X�q��D�4�:�g.���W��:X��A(?
���Gj1RI�I�?27�X�5�����l䵮���׺u���
%@æ�X~�윮� 
�v���q`�/5;7�l�Ua�1�/��2h1q��$=�nփ	mUz��������H���ҷ݉B�oع �. K7�BN�ka�S(&�<@JA�x�K9?,������e$��4�_+7�aHB��$�K����"�����"9�*B���_����JEYK��*�i�nM,Ad�	1��������Ǩ����85�`eY5�%����rXP�RI��g�",ӊҮ��@?����A%��(.�z�ӫ�=A@��^��	�6����%��rҗ'ʬ�+/�96�=i�mL��5G��-G^�3��I=��/=�H������޿FY�>�KnD��5�	א�{nX��1I�o��.��Df�f�������:�%��Sbp��bZ���CQƅ��,���ԡ�=���n,�,�}$��I�Q:��>���?.�3��D틯��_�%|P�-O��MH�;���x������� �� ����`8Q$V'�M�W�y�ߵ�/�F�B^noQpS6vܷ��t��2&Ʒ���M��&jVo).�OVB2�F渺 1!&L˹�J���� �������_U�x���!:�+'�Gd����6<��D^B�~ߤ���	c���v~. �~�ٰPc��!X��Y2��hn�M�T�K,�� �q�Raֺ�z�
��Ƹ\�}֊�o�{;���{�|o�m�Q�2r��|B����kp	`�	M|c��ֳ��U�V9�@��$��c��@V2��yۇ�I������B0��\:n��)x�	�(~(�R�y
5���|�$�s��F𥍡���Y-|w�6��*(�d6g�X�ַ���f�*�����JW�qr�H0	��j���NJb�	t��s"5D�
X��ײ�-�oE��q�F>�P�\Ǹ�;t���I)�=�����d!-L�7�e���.�;�m[�/��Z2�����lw7���;�%�������{�*8�aW�d��i�`#����=U�E\U!ӥ��	DFmi�����
|��F���5���:xč�k��=�X����`�y4���gR�r$��uRjfKGc���Oxg��*ʋ��8�)���8j_�e��^�1����2���Rx&$�T=�pm[���e�0L<$��2������<V2�r���Հ���t�� d��.stW����Z�	qN\i�1&pZ�����e˸}I	#�g� o��^�6@����H�r��Q�Y�ݯ6�p�k�@�W����9L]wa`��܊�[�r�M�ӿ���N��:�I8��K��"�+΄h�<��o9�->cf݃�� n��|d�'C�!�Q��J+�<�Nu�5�(�^����]z�1�������$|	X�L��0.Ni_) �۫��5��7#5�@����t6x%خk�x��=���J���Ea̅p���M}r�G����%t��5���ͺ��SNA~�����������EB�t�����T��NAx�}���|�6��Ў�%��$b���ȃ�+E_G�ޥ嫌�͏_���v�N�1��4��i6���#��̶� ;5g�}o�:��KX_X�$c���;-J�}�O�p�D��<!+����&_U �xu.���P�t�5�i�v�_�)�����i�ۅ�C�ERm�ďcF6�7����N#~4���%Ah*	m�S�ƓrWt����q�Ld��) *���ܼm�2MB��k��kԬ�ϞQ��La�<z����� ���\���t�l�h?0�Ke�c'(2=e%�:S���z}Ծ�Z����4oS+���<�\ܥn�g~���Q�VTǋ��b�K�=� T�^�h玞e{� �]��ZJ�3������U��t�0� ��a�Br����
m*[,����:X봬OQ�Jc ��\lxo%�l")��)KTb(_S���!�~)Ym��+��)p��Ż������?����ڞ��]%2&,o('��7�9<������7
���;�	i�9G2@xVȘO-
�Q~J�j�a-I2��o��e\��x�Z�ETD��L�E�H�ѝ+:��S�.���K�N���;"�Ǚ��1I���`8����g/{|O��'�B��Y ��ب>ݽ7�t�ǉ��nR��mǋ��ISf��3��L<��0�|�]�1]6�����$Y2N�x��p;�|�@��R��o<֓{�;�ͭNHv�M3%(�B=��Vc?�[�{ ��	գ?ns~L��������� ��R.c�� \O�u�J�e�:/��_5k�Ҍ�āa~_����=�@�j"��,����P-Y(LQ[�͈���^��S��'���l�����7M��:T-�W��F��T�DM�7�@Y%�7�@�z�v��r�NO5�Z9�1�� �Fk�p� v�Ho�y�0J��y��Ҍ���U�&��3g���ˌ���s��h�D�j]2�	KRԳ_b�k~�����z�
-�M�A�7y��k�ַd���`s(���X�=������Jw`�h�8��ef��s�g��<�r�5S�Â6P��%r��}�XF�aI�����ו��P��j���<�����L>}�.yW"]`��JvJ�b 빰cI�Q�A�wYϟ�"�����]]�P=ja��tm�ћ�c�U>�#U"�2Ň�7 �4��f#�p����)֣[٤D�弓����ׁ�+�\��wI����o��r�q��Z���&�X�Y� j ��y�J�A�P/7Yp�2X*�N�|%Ps���5�[㩔o+���\޸�J��v	?�����9'X�����t(#�6���>7M�;��AFpOrK��	������Y�Q����+Ι��ơsR�ݑ��O��i�M��u����3'A�1il��M8fM^��	�����������G�X��o�y�0�}fm,�����Aj����ly��`y�o&����c6�@¸��ay�L����M��C� �����&��P�`Ѣ�� +<U����nx�2�S?��܍*�<�<sa�1�΀$~�uz�I�*�������}yǞ�.5e#$-���l1%)�_�U�i��*��o�N�.vG����ّR��Ȭ)|/b������ ����|Z�-�y�XtO�d:�k�
78d��X& �"��ȯ=��FE}gꔿ�7Y�1pf�饕�Y,���Y��Z^Gr�q��r�s�]{��Pkh���w�G�}�ûC�ɽ'��Fi7���~����6Ub�d1��e�@�'!���n�Q3�ؖt�W�r~/�K��%Z�ޯ�l��?Y�̎X<khh`8:��C�bp�٦n\�:�~/c�۔2�,�f�6Ɓ���\��SHo@���8�����Y��J�9�[���`f�t�f��ϓ �+&����l��}#���ܓFT�@��6Y���l+E���e�o��t7���a�0n?t���G�o��X�ҧW�W��;�A� �%�o�����W/�
���e�I_�*�n#^G�%
?�,��cB[cHp�D�������p� �g4��<0�/aP�Q#c�*+�[�=C-ۍ�T�v*Us��HS�X��`a��BrJ��uV\�������H���c\��j0�ÝV	_!  %���]������?	�Z��T�z�%"!x"ʺ�=��!�)��2[�����?�h�n/[�QӉF+n��*�?����һ%R1d �+�D���?}���]�C��kE"~6uk�5yJ��"�׳F�����*m�=Q�y��Vb`���BO��}��EZL����\F�C"%�T�GY�^Xuή��&�M�����=w��%��m�W��{4�YzqP"��ė(�8aY3=ˍ�Zw~�װI�-����ϻ�u
���n�&<��4b�5��	M�q�+�Ӿ�:K9���C��7!�[�j��+�@&���qBW��o̬L��5#n�1�Ⱥpg�Ɏ��F��)9��[�Χ�m������C��j��Tx!�D�Ρ
쌐/:��J����<�˃L5��	����r�k�^�9�Ȍ�V��3���H&!H!{�����?5_�K>n^�#�����]!��-�5�X���*� I�A�7\��I���[=�GŦYl�61<�3�6�O�=L�4�2�1�Ĭ�0��D[���z�F��
4��6O�>̌�$��%؄�P�6�>�?�/R���Q�q�g�Vִ�yYv�cgN� ����6�����n}�)�Z^)A�V�e�@^��ı����P��G���Ku.j��Zu�� �0�����4�VvXlxV64EB    fa00    2bd0&_L84���e� �M�������g���!�in���|Hy �>��]��`@,�v��$��V�	
�s�`�E�I;j �w�F�a�Ȇae�{�m�6���j��P�'�\l�mt��&6Gx��&`�����qQ�9�,ʱԛBȇ�b���!��w<��_k�o�2�qL�<���=G_3�����F��LN3�w�*Sy�K�y�	�x�&���j��7*z!��]��l����#4���ѝ�5(�|�9G�Cͮ:��|�	��5p�õ|�!G0�8�Z�A��٤�j\�&��x�]|yk#t��2 ��T7ǎ>���Y�~�q5�v�Zڱ������!jw|M�p��I3��� �8�
�zR���_t�����|���)u�:�sE��xOhfD��)s�
��㷸��]�
҆��>�㦡s`��E(s����<)L���m߽=�!�0$�#S��
b�>~��w�ba����p��'���z09��
����o�4ק�_�0�h�f�+Z��upۓ�P�C��U�������3��H��֡���ben)/��xL�N$7�6/�r��a�]�'�g�g�=�.����'���/�X� Hf}�D�wUy�h#h?	�:F��+�RRuE�ofPNn���{�ɈMr�9�HW6� "�=�{�H$KB�e(�RW7�n�曏(�������b���l���eæ��Z���Ȥ�	�!� ��K4�$���{(�&o,[z���)ܱh�D�P�	���p��J��EfAa�q{4O��ʃkpoh�ܟ�8��#D�9��y>a�Ƹݪ��/�~����@EW�W�����f��<.����)�^���W#;Ph�`�N��Y��D�ai�F�t�O6>%o�S����s��r'�d"*�,s^Q{5�GH��}�[�9䄵r�L<�H��z7���"],�ҋH��]l��`��S�5~c1�ߣ��{5��ye�9�:�j�W��m�1�+U/j�4šsd�o���	��1�"O} ��V$���[O� x?��Ċ��f 9��[7�����;@���6��ˎ{e���^4��J�o�iU�w�b���7�1"����HU A`|���!�>�������JR���"�0��,��ۓ��E��1hH2_���y�~�A5� ��^e �aR�:R&�?/ �����q^$�Z �BpLό@z��R40޹
E#��� �̐�|�_����SK�Y��Kk ��0aJ5�WE�LR���7����{���'�%�@ωq��i��s	s�ǥ4�#4K�X������@��n{ �Sg88uA���[���4����M�U���e��]������]��F�"�#����|�3`l ����6_��,T����"HU,��?��;p��s�u-�`�1����:��v���si۴>�D�%�L�I���z�q6!�Ř9����8z�df6��i��KI���MsLr����%���7��乩�)�����|t�&P^,�:5Q)b���b��$3^���g�`3���^{ q*"�2�˜��i*�E�i�`�L��ʲt78���K��L���y�qm����JR�w�����5ҀT����U8�����Mf��Y���h�y3R�W3UxUe�BS�J6��h��,I�5�T���r�Q�����@ !�������KP���S�J!�2��r�&��s�yl��U|�V�j���}]�%4�Ǎ�z���������1�T
߀�0+�8Z@uY�ߍ$XG���!��Bn1o}��9.҂�<�m�7S�20�7�����h|$�ߩ��A֋.�;���K[xZ�ėq	����KԆ�`q��,I��;I��q��2�H��yRU�)�B���d���P�����r��af�2�z�GA�+%�vf\QD_2� �c�j,t�u8�����H}t��2_ǰ�ڨ��s`�4)h�j�JL��zK�fm�H����5�s7�+���T�=�\%IC����x�m������Gp��:m�x�FW.�P������Q�H2����� 꽂�6w���dJ�B՝豁������ZL���p8gn�3�+��W��wP��1O�Y.�IeARokL���q� �|/U���36��ה�n�+�oI���|J��
���g�u�M�U�����_�;�uX�h��*L�=��&;Qâ�z'� 3���_9f���Ҋ^�|�p
��%�G�zQ�E5�2۾<D�)�y"g?r�4ޥW
�C���}���DnY.�6Vv�h�(a�R��0�.����T�N�d��I��٥�Ie�\Z����ѨX�F;A���U�w@�D��(��~�� ��8K�&G�=N�s�ܯ�NS֥�c~�B�g���$V��|�FIH-1�!vU���t5�nt,G����X1��x���o�+0����ؚ���5͵�"j3h�`� ���!�3TP���^a$7�Y@�ё����D��l��5nW{��~����[5���R���}�����t�dKj���]P�H����Ȧ܈w�80=�R��2�%,fH���2���pˬM[��M�7W����/c���m�l�)$x�����w�.t6����@��^jݶ_�Kb�����=h`��
)��;/�9�r�LŜ��7��:K˸E�l�
����3F�"�����yn7*aF��ZER��������ĭ.A�w���_j��5�ޯ�.��n q��X��Cp��ݫ�
69���So}���3+Q�)B�/\�~i��]���x���w�.i��| 6���ᡄ���Kk�s�G�_�m�4j�H����6��40n O�h���S��zc�Ki:�
���h
yۡ�d�R�VQ�X�T��1���,.�ڙWݵ�H�{�Vc����f���ms��M'�0$FߢW�� :�uv��J���\N�?�l�Q�mys~���ݽ(�9iCb����?Q�)�#ap"���3լ{6����mv�K��fb�b��i9w&��W{����juL�VY������[ur��J��WnjtWR['	.%�Vh_���l��1�P�s����>j�ў��m��g�4H>KO*sw?��X4��O4��e�);���J溏waݮ���S�:� f�2�g�Ug\=	i�.��0��g�D� 9�Uk/���������_~��S�CPY�FSD)���ݚ�dLO}j��[L������.��*�����k��@��v)9�d�B����i3W��
QwS{��hQ���Wˆ�b֨{��K|Á{ֽ?G�]Z;¸��NJ�������r"�f�k����b�ߪn�(����ѧ^th�eh��j^�9���ɜK��l`}�H��"cyI�Ȣ�w
Wi�'\i+^��ōZ�|�)	����r�0+�3����|�% ��7^��2�P�N�ӻJ���a[�<���閷$O�*��\ҵr5l\=Eܝ�:۾�,��̳S�s�Y�	��vͿ*��:�*nC�ޝkjR.��?����z��`@���4��v�y,B���+��<�Y�!Xr�a:)RL���;����#�r�^�{P�`2F���T�cMf�{�\��Ѐ�M.���m�߯�/�R{w���y�U)	�1��@�����o�Cw~mf9Xu�N�Ej�+�����v�U��L�)ۃ�-q[t���M��@׌��~:q��O=����Q>�?̪�4�w6(*-�%�,
���h��r~�i�� �t�U]990"�@E
*~�t	�8S�l=�r�~�Ge4��l�Ȗ�[�/)����-�.��c���0�M^Vx?o,�z��I��Dd%lΟL�!H,d��+���7�4Z[�8�����\�Z���-&>�7[7�e<���-�A[:fb�'�_��ǻ��7�2�]
�,3ߧ�lEw��e���!�����Q��]GC����u�%ikhgsjHCˢ�S��� ���Oa��H�`g�~V��`t+Lo�w ^��iΦ$�X="ȅ����Ҙ
��t�R�+\,�L�_����	�| <ס�6��D/���	&W�i��y�,-��Y;�k8K	i�J��x}*Rz���0�~����yYF~v�M�Jb���蚢�Z8y��7 S���s��m˃��ɦ0�~ޫ.pb~��4������w���z���,,n�Egj�w󈌿4.sݔ<-0/�^3�}��qi�-w�z�Af{
��y��޳��:ݶ(R	R\����,�Y��;�B�E8v%͑�=�0;Ȍ����h���t���%E���Nv�u$�Hw�(�?���b�Y
�h���܄�d��1$��Ip��ꖚ �9���(+O������T[�X���N�s� �O������_<���vd4	6�/���9)���d/'ӏ�y�SW\Ny%6��1]���vw6��؉cn0(�e*�9J`Ӈ�p̅��9Pv��Րs�+��x߯��cJ&�n��r�a�kŤ>���S��S�/�/v�8��
ԫ�8~gC�ļB8��
�zg{���r�A�Y�.	�]gW��H��ksܵ� l�1�����Y�[��X�f#nF�w��?��������Fd�_E��E�S��Tx��TJ��.��#P-�"���X��'*��fN���I.<l�������8"�Y����ܮy�(|b%��vy=X�A���˩@��xm�Yh�m_P�������;���Ս��*}]�q\]�k�9�����p���5�|�K�3hN� nɩ�@L�����h],�"]�F���f���zuF�눁s�"���kVF�\�g�C�x���d�x�/g��p�����'�;"��ؑ]jSb��[bTq�g���-ܲ�[m�S2AK�ݰu��"FG�����ۉ���;%G&AU��DoӜMTѪC�U�3�c�$D�����˽��+����]�=�~C] �B�#vm�e����c��T?��>C�K��l ����7z�A<Qj�Ύ��V��@�"�{���S,խ���2I-E/�,x(K��P�����g�l��.�k(��ɱ��\q���Io>R9�g�az>�3Y�^�D´�YI��
#��A�+�/AZ�q���#ʬH��Y`v�ChV��	�f�ĵ��R4x���M3i���ރrnKu�	�x�L��_���e����0��Оqw/J#���'���[�[�Ũ.�i���.U5$q��b�}v�[T���0�t��5�o�O �[����Nۙ?F?�y�����'��	:O�pMΝY���6�F�[5i
��u���S��jc�zO;������y"h8�h���������94����?6-9L���C�jҥ�8җ�Cd�Qd�4Ї��l+l|�5�z�$!�m,^hT���S�����ֳ�e&sP�3�1�	��ʮ���J紕�{͝WYf=sȉ��|���5��l�=�� ��OϾq�=������V�.��J'넦���kG�~��E���b���rm���Y?(�=�s0�2gR�54�@�Q�J\Jw4�l��ң��U6�6��`jMTOU؛h�Ŕ�cÅ������ً���>
L9���w���#Wd�<��VfK~,�:��x:��Hga �UA}q=�H&f%%򩯫=o�'���6���Em�1�4g��x2b]�T��BpLS6|��#�k�Tp_�Jj��+W;
(}�p�Z���MPx�4`���>㭠:�`%���~ƾ{q�f��T���k��_ʢ�ֵĻ��N�Y7Yм��0�����W�
p�v:�`1fK N�ҕf#H tGa�KG�7���2F�==�U0 ���p~�!�$����~�a֞{M8�DOF��>/��,Y���9B����ڽ�kh��OOY���Ѐ\��d%+�FJ�)\o�@�_����ey�EF����hu��`Ε׳j��'3�t�q?Y�os�_x��,\�,�ܾi�7�ش-	t�/WM4�3��NZi���%]�c­� ���k�07����W)���PF�<��֩�]y��K��B]��\У�mha���^&��z�1�\9s�R�~�,1nx���J�pe9N�K�����3��j�W&��}#��W�N�`SJg^\���s[�ʎ@-Ƙ������b�	)qP���g`</��ͤ$<��?����3�..v.:��gR,��.3n����0�wK�.Mw��E/�c�\Ĝ�=�ם�$=��ja�uH��8���O��9����<(\��k��60�g�*2�������SE}q��wQ2*��һ�k�ï⼘�,����ˏ�s��O/���t�2r�?$��^��{ >�����K���49�E���-��=U#�0Aޣ��>�L�FwL�w�\l�b�%�
W�g�"���ӌ�F����p�5f{���DS0*�
��Ղ�;p��_�p�p�of�����4��}�}-�E��v������� �皦��[���ܗ�3�?���
��\w]y;��UG���#`�2�P9Z���
z�W�q�}[�kʣ�ұ�zm�P�C��K���0��6��c��/n�_+F5}A�qǵ��et\/Ӂ�l���uX%P�f_��B�/�9g�ܯ,{"�v���{]±mJ;�Fa�ɹ���D��a=���@�ͥ���
r'6�|�܃��37�P�����e�7?ӲF[+���2)�):���U�_���q0�~)�b�(?�i^|R1Wg��@L�G�{��B7�0nm��дI�+P\��&Ӵ��5�O�l���5����9�������k6\��-��"'�3X����9W�|=Ь�z��$�V�m?9u<��R?@y^����t�SI���<��B`��ےP]�Ǭ������,�);W�=�8��&�\�@&K�&�=�*�����!ay*��-Ļ��c���%�TCz�y������B�%`z��_�V�.���u�y/=��\S~N�5
o�V�'��+n�_>�聓�� ��m�-����PE� �Xn��������\��i#M�wQS,X�<-@�h��<ۊ�Ȣb�:1��b}�E�����l6 �U��5
����(d��!�+y`�<51V�j����ֶ<A�l��*"��rP:3�)�ZXʍ�Y�xݜ�}7���O��W�	I��pN���8X��r?���t����Q�hSʰ:�}g�����)��^T��V6������x5�T{�S�����ߒ��Z���Vr�ٙ�k�˴HUPq���~�3��hs��ͻ������+�ɂ���ǻ�@�L/�"Ӆ�����H8r��I�Dދ��V��Ƅ�G mOH27X�,�p�� �[����۬y8x�#aD%Id����?��\�
b���9�c��Mq�,Ϛh]9$fY�.E�Ҷ5��6��H�6�|��,�k�q�Wf-�<խ�*j�#FP�,���ǒ�X��6���!�����7���SE����ϝ�D:-k:/`�I� ��4�� �s&"�Ͼ�+R��o3H*�$}���M�B��Y�C�Kc-/&\��c탒=��\���`Ҍ��5]��K�Ҝ%Uta`��5.��l�{��X�!�?O:g�o��3��w8c�_�;�S)�tQ�a���8r����c��+�����6��J�N�����å������{f0t����+��L�qʦ����=
�b�'%�ߍϱ	��4�Γ��4�y�B�K�<��7-\�uy����	���A�_hd��HTutR�;��O�tq���B �>�6�0�w}�ALj�D��s
��/B-.��
�)!%����H����̀����c'���/PԬBr��MD�p���P�����%b��9�y!���m�����C'��ޕu�U�|��1��k�z@H��{�(d�_��Gm)�<�T3�ɕ��	Z���<A�2�7��� ����b������p���}����^F���tv��!��Zؓ���$M}�/����."N�ܯ���2�6��Y�8zjv�q�y:��g�X��k�GkÅT�LA=��/V��w����R�$;~F�yv�)"��pw���^X<b	�ޣle����7�8΢M�{C���!nd����~�ـCD��l��.9DVJ���ж+�
vǐ�(��{'����93/؋\
��D�����{V-��i7����õ�mgr<�K�gJ9m{������jxK��4�
�\�D�*HGJ�uH����N��Ж�RQtݛ�� ����7Oڷ:��+�jU�b8���jp6���u�e�d��p�vO�-�/�}ש�F�o�g+B����8��Q1�"R��e?������7����B����dH}X�K���hG�+Dl�B��"q�mՅ|+�A{�_�6�'�m����K���%���b�?�]�E��r�W1s��h,��Y��,DT��L\������_]�W^�Pg#0�����mn������d��-ڋ�uc&]�KC)�&��hc.���l�2���̓Ս�n^^�8�������R<U�sR[�d����q{h#*e:W�JTGѸ\d=o��[0�-��Hn�t퇸	�J���9-��V��ϔ���~�ИPG!����ޣ+����ɷ�{a =����Lw0f�U��} Pb	1�m�EI��	��SX��'�{0�8�H{8�v�R���	��$��wi���m�t�	���+��g�N�dTD3#j�����c��TjM�t�v6�2�@�2�T��bt�c��Ea ߻�E����sn]���Р���#���s�^��Yax�;L�95���)�4��6z�/�2���z��CF_���
�q&��Hu�ţ�$�7�͋K���ϥ`+�y���%�s}�2,�1���l�?��'�2��d�h�Y$,V��Y.�nf�����2���"�H'&�jl{|�����7����T��]�<p*Q�}<2e4-�ri��5��s �V���}d<ޗXT��� H�^�~���5 r����"�Mу�v�^����+V(i�㜻ި�	;VG�T'��@(1l��DB�k��7W�1f
�5����9�>�c�4��ӫ|:�|h�x��X�fX�����\��&���	��ΰ`�>�=CL�5�QZs��h��ϣ�\b�b��p��*^�Ku��i1G�z�̝��9#F֐��wli�_l�*�P+~�h�ܨ(rb��."Z���qM�Uܒ�R81 �3�sߖ%H�r�&�L�Be�֘�h4�*�7r�1�[C}�Y��i@Y�Y�#�/F6MZ��vqQ�l(�1�M�AD�b�T�p��ꊄ��d��r)�~v>���[,��ǩ�uTNMhF��Z�����hљp7�T��k+S	#���l��<���y�D&���e�U 8��kOj��e�OE��M���|���8*�Ÿ�0����~3��6���/�)q=O>xӴ߱NN<%,܅�r���, wmY��5JIqv�X��u���_e�G��N[|8\�O�	���1�R���������MܯG\ʽ���%�������<پ��R��6f/��3OH�h+N�<a���K������p���Mt�������l����u���,%�=���I�s�3�Z�;��_�i�&�F��q_i��*S�����<(�Mv���8��Գt�;� �C�(uF�l����̆�9{P��|i*�T�| �d N�������O/���B`s��5׋wU����h�q��W|BS�äA"/?�������K.�2����^\zݛ�^��WV����Z�����):,R���-��s�EVY��*2տF�ʬ�f�kE���r����41c5���I���6����U�x0��cG��¬\b���u���6@�iҐ�Y��P$�eԗ@�3c4�,�Ώ��]&��3�*���~G�t+�k �Hs�3��t!I�/�����i�"�◄P�"5�A��/��ˣb�LN�73��G �q���L<cD��*�Б�`h����s:$�kঽ`um�B�m5��s�^����z5v�yD��G�{�0½+.�)�I
�BB	��NO�jO�v���ѡU6�
:���z[xN7��p.ңG�,���V����G�.�v�gCR�ۉ{T2U$�+K���G�LC{�B��L��kq/�����}�e'��}���~�ֵ@7�Жd����ף��̓�+�ƭ�E���+�\Z�������&zc��YW����Q`X�҅ǖ������c8�C�T�gi��׈m�p��E^*�����{�p��̆B- ����z�3v>��u��Ž�G���A[��DL����^�rIi����T��}�CN����/���ͷt�9/t�W�d�a�[�1$�V#���y�l�L�}�%(^����a�n��M��E\��- �������Z��5�Uy���pR�v�
}���QI z��?�C�6@i�U����>>aq�u0�.�+�i=�����f��pm��v���(��G��χ@�,Er�����#'' �JH		�./��].�uhz�?!����e�����[}�i�n�����C�1�� R���"���E��Ǵ�"b[�u�>�{߻��>�}�:lK�RT���8�G�0��LDH�*�U�vD��*���Iئ�v��N5�����(a�=���J 6�Ǐ]P��k�>~8�d=p��/k<�[��֤����E�N�O�ο�4/-�*b�Xy�N�Lj^*KD���c�%�g��(�j��1�K��8ٱ"wv]���ג�^[u4�ҍ D�J��rDL�,�����M��/�9�Qs��3ƾ�ý���<=�6e�a�Mp�	��z�c�
����lK�>����n�Z*U�y~�qr�!��b<\X�S���4Cد�q�A��|�X5�ՙe��
v��~������F�U�;�}D��ى�2�f���m@�������-�pW��V�~;�ɂ�m�ٹ���;K���T�h-��j��<�w�.ϰ��wi�V˛"�)�v��_��^�u߬0�@sz����T��E�>k�/C��!��qwg�Υ�U$�t"qa������XlxV64EB    fa00    29b0��{Ua�2�V���;�DNt#���ˠ�����Y&�$I��(8�5^A���+ګ7�R�n�����z�0Zzp\3��p�XIO����&ۭ $A�8EǏm�M*ۅb�K����z�D�H�����i9r�G�È:8��F����f��:�����_\޳^�<3��j{Z�hW�@���Lb_�"��-��1��Tդ��,�`�2��9�E'b^}ͳ�^�b(�m�:���J�>`9I;��wt7�:��J�	�
��̿3�NN�\R8�>��a�l��
2}�𶼃���kN�̙�\���0f��s!v�O׷���HFQP�	;䍳@��h�,���&�1�y%M��~�w��P�K�8�Y�3�_{��ج��nI�PStDN��%�<E?vG��[D��/��5�ܰ�I���tǘq�5i|x�o
?'�6E��N)�.� �Yg=��f!W��:�\Z�*)ึ�y����[�Z��:�Î�К`��:�z������M�6�V=��.P1q��6������e�o/5i!c����>�u�``���z���y��x��"��K����_��b<�_M<5s>?����#Û9��$�㞌c苌���BaqE%���c|�	�<���T�C�z�,^�3'G�&w}�]]$_��i�#�������=���Y7<��f��`Uʆ��3��a@z��)������!�3�x�l��u�k�o�&j���\�t�SO���Y�r��2覎�{�	>���); �e~�+)7^�r)-x)�X-�B�"#A��iz<�v�#�:PgS��P�"��˩�?I1ߣ �W���av��&]ǹ�m��j1�U�́��X֮*a`sɫЌD���>Rc"o؛l��$5yku&���P ���ZV�����W8�i,�8��;�q_'�o���97��`࿕H8ms�1O�t� ��c5��0x�[��֐v��@������~����C�PյN|��5'y��i�y�Cc��c��Y����'[iU.�	_߁��}��C�>��[t��"���9օ�׺u<���7�Sv81L��i�6$"��	�I��,�N�(����+�B"���6�!�_�.�������¦�R6&�ג�s�6s��� [ݚ�^띝̽a,!��T�D@|���D*�����Q�Yjz˘l^�h����+5�"ʊ����{.��le&�N���x�s�,�g�g�Tl<�ek����J�0lћI-E�(F ߏ���y`{TG�6�k0X�˽�0��=:X5�Kԇd:Y��Լ�	*�l�v�q��c�M�U���:ة��t�C ��念�#0[���8��J�{4JoE�X]"q���\"<.9�ch�?u������m�wQS����4ƻ�����=�m�b`P](Wtǰ}�b~�Js�Ͻl�"���=���_O&�Wf��#����h��n���l�U���͉�",�N��I�8�w�?����>�ǡT��E�U
������
�P{	��E���,��Co�"�>Nc駊y~���搘�VA�e�:5~Q�ް��E~�4Ұ��GS���P�%ՠ��T���J��cYe��
����0$���]?��~���+$9h�2��G=5��z*"�yŅm��fE��Jͪ�r���GIq}�m-�������8K��������U[Ǣ0�&#X�H!m����7�y�g�U/Y�-����U�l���}Z�J�.��煋6���h��Ƶ��g��Dm�Y �+�����H���F�����s�
83Wb�8�6����"����6�fQ��	{*��w��f�[B�>a��ՠ���������.�]"5�b���H�Q�	�o� ��a�V"*Y����*'r����|�Ż�FbV'R9ב�n��*������������},�[����4¶=�8X�dD�Z�EX�ލ[���k-��4N�� �¤����A��R�c'fh�ʆ̲�77oL��!��x�6\P?g2�I����=�s�J1�A$k�e���W���m&mt{},ճ@�YC֚��ĵKدO��V�=�}�$W8�;��Z�N�� +7<*�)0;���c-���G!$�$h�XOp&�3�o^f�}lG<��c�O���IC�'ء4-��!a9��ٽ�����3�_:H^��sΎr*��G�8Ě�7~���
i\���8�� ����%� �qW/�By�K�ޣ��KdUB{Qk�S�]�ZWե��w��8k?.�T���,+��i�(�~zc`��Ժ`��T_�u��B�n��ai}��!Ճ�b�e� �	��(rw���hA����>��7�ٓ����(� ���+~��YDqc�6f��W�����~~#�}U��= 
�f�1�+hf�������5�à�0�N�N.���d�Y~�fx��r&���.W�/�G�c��Aw�e����xo�kI4�9��]�e5:.P_[�e'̉�����~ɘF%Oʆ(R�G-(��P��z۽< q��Xk!�^��*E>o��1�%�����\Ff��f��;�V�c��4��C�p	����^Q)��	�:珁�PEIQ�JXp�c��W�ջb� ��L��8�qW&�?6���$D�곂�`�P�� �2�Ŧ�3[���_F/�ą:#��$V���E�^�G�H+����|�9�� HG�;G�4��3�P׍�^�Rm;��T���ދ���M����=����t�?����"�C�{�M�k:`��ӥɴi�d�;���,��Lb�N����i}��K�ZJ��sزeUR���B�ϴ	�@աi�$92�ypfz={��e�9c�eZU
��/��,{]3c��&wf��w���s����4�cDۺ��F��q��|P���H��i�+��¤�\���G|�(>����f�R�S':0]K�����9�Hy��E+���Ŀ���r�Nؔ6�*fuYn��~��i�$�ٝQV��kE�J�%6�1%�YU
}U�`O@�|X���Nk��u^7R�:x���PF4Ðz�}���5�.�0���0�O�ҏ01�|��a�0K�$�B`�\-߼a�&R��y�#>n_'�N��_�Dhq�����h�Fڤ�Ql�.\��?5S�� O��Y��A2�O�t|�؜���%�xj�H����ø)vs��J��{��9v�v�V�?�B4c)O��n�mUC(�KB��P���q��\T\�a��܌' Ճ�X7�N�$�u�ʦ�3���4o>Q�V�t��FO��P ډڈ[�_�6��l��"h�R�O6^BM��9�M�f��!�y1E��t�0X{DaV[���C�QH3z)������ N5�����N��R�^R[�����7�����E�bE]�h/�C�%Ë�<Gґ��%�d��ƣR2�;���Kc� >Y�.q��5?�S`�̏�\�q_p��"<1ev4~;ﾘ'�g�쫐��Qz}���G�2��L�/��!��Y#���57V����L��`(���2�:��:ĲN��<]�M���cvV��dPЂ�P��ӏ��7�,̄Mn+�dˇ+.�Jaq����岞�x��U>�^��eg�V7�bߐ?f��S������W\���F�u_���
{�du!s����e�R���2? ��8�B6�].����o�?�É����e�r���V,/�m���7���B��D�|���Q�In������	�Q1{�������NJN�#���S����+���ŔLDV����Ĺ�ҷ��:�}�p��F�jCi!Y~`���z���Y�����[�Y
+ԫH�OX���� �j;��<�J����SK�4#�� n�-�ԓ\����%:���ߨ��.|�{��M� �>JY���yw_m�|'�[&r�� �a/��
��'��3����
��脁�^�/@vać�I�.A6,�TV=d���q{��J�^bg QWz��mi$�}>e�y\r�ս��D�M�D@�JߤgZ��
�/]L)�)cT.~��A���w���%�i�g]��J�y�Ȼ}��kt�wsLh�Uv�!���������ݏ��.`�ZE��QIW5����4�	ￍ���g��w�B����Aj(;�l��<�N�q�N��%E*Dl���	��^�w6v+�^T���j�-���0�c���P:�}�����N�[�F*ꇜo�� ���dkx�=_0dn�J%�B�Gc1�Bä�U8�ס�ٷ����po|�F��&.-�˯�tt�nD
s�R+AdQ�	�h�HPn��#�^���.Y�J2�D��� ��Z/z!��"�6ZBh�O��U�RP�"pO.X���!�����?����xt9����5kQo��x�G��X�Z0%)��;2FS����rh"�}���'���YNÔ��*��@�Zn'��A�5�4}=��gy����ax�ż���8]����� =��t��,g�/��wzo<5ɞ��/�6[rЉC�c�[>��G��\`���j8� ���� c,.1�bM0�l[���]�z�j�8��=(s'����qsH�)�mZ�3���c@�(�YR}^�/3�]Վ������D���X��A���g�
0ŉ��-�������'��.+<�3-ߙ�����yK�X�p�N�X��!��U�.�>���{��=':X�]CB�EyJ�Fc�b��ᚚ�YՎNX�PQzΡ1��*��$Of���ئ����U)����!���@܆"�/h؈��[G��̘>S�{7�Y�̆*,*��o�=���Z�ݻG4ٴ��b�4֜P_�@Ff���;�ͮ��S�2h8Ϸ����rih�Џ����mVM��8���K��t����ˑ����Z+\
�u�X���9���@�tG٤rea7١t�|뮛/�Ni��:�c��b|@�^�0>��͂�N�V'����_�����e���2�{����x?��,�H�죁�HÊ��Z'�M�E��:�X�Cb�)>��VP�d����x(��w �)�X�S0����5��G㚭I���ٮ>�d�ҷ�\Lɚ\Kc���Z������GC�%�8��XM��KZ5f�%�)h������#k�4�r�q�}�N@�e��ِ�zd��fH�!�{T�^Z��c�oip�E�
��/P!���wh�g�vΆ�-B��֒�֧r@�&�}HuV���m	+�*Ld��8]Œ��EԜ��!�6`���q�jm�D\<��ًt���_�%��Cld�aCS��nͽz;��"�C|���M�=�EP�2�8#�lT[i����$���v�4s8��������ڋڿ�X�z�� 4��ʞ�U������b�� xb>�=�y7�.�R�5�h�!g�� Ε�PM���-���|���b�k������Z &]ie�4û0�<2��!˼�Fuo�kHg;������r��Jvvsvh�jGQt'd����/\��]
��V�I�F�6�e4͔��q��g��~v��On��L����i (�ciu!�v��N���ߒ"󢓁h�6%x��@~�ت�����
��H)?��2}���lYq8��_oq9:�?mf�:�(�3���!~*7��$.h���Zͱ�w&��v��/�3�Ww6#�o2���P6x���#jOS(2�Os�t^�Tz���%�Is� �S�YN���Ǉ�%��\2z�=,��IE~!��t�u��/rvm��]����?* �M��\�ޣ���P���^���48��jTAv�������;~C�E�X<��aF�4)"�D�;_���G��Q͙1�HX�&���K74�,{���ޡ�/�KK��J�x��S�/tq#3�n�ແ�Ե���	8��r��p_� V��PmΤ[���|�p�ϼ��g�{���]�8cҏZ%Ơ�#�Ổk�*�7Wߣ��ߛ��Ћ]TRP�^]_4���1_@���x����ޙc6��JǧY�{��I3�i�.�B8�ye��-�b^��.�ZK�J���"wv��ܥ:R}��&8���̑)�ظL�6�������!��΀+6@'�y�u8�������l��JС�z��7贽^�,�um�+0�;�֠�5���py��ߕ��c(0��)bi\aaQm%��E۹
\��e�&�M#$hɉ�kgZ�Gʟ��މ�j6�͉K��m�Ϣ�cO�f�_K�6��\��37 h�-��L6�
�*����	�~}\J'Ղ~��Gn@�$DJ���S�xs��������Jߘ�s">8���'�e]й�H����\�X9���:B(Q�D&	�B���\��Kr����<�g|�Qt��pc�@�&�_p׭��;���y���jv8�Dr�9�!N��z��n6����2�u����d,Oz��G���F+M
��?���\`V�q�B���"c��t&'<�ՠ�#���}X���������p?�7��@��m5@NBS�O?���/P�J�Z<%B%W�b�5��
9$��f|�V�+�P���䛧6w8B�˪�n�V�O:zxV�x�v�yÁ��7]ً{s+�DH��2U6��1c�p��l�d%v��d�����{/����wtd0z�I�k���U�H_�Ԙ����"�_�R�7��Q$�vh���l�>4�����^nnl�K#��N�Wn�g!=B������Þ��HC*�gh��N����ZN���{	�,�@̙ߡ���{#b�ְ*�g͏ڼ�!0.���yfk�H���M9������ׂk� y;�o�_b���Lu�����歔�� �*yinV��O�M���r�`Aՙ��kD���ծ��٪�6�����f��7��:�$b�
�V���N�"�����#�@r_��C��W�����М��?�?��;�tըH�?F�&�g��f:�����1���Y>z�;�\��?�:ٕ㽰L��4�D���_e\w>@A����5�xs�-�_7d|�YI���+��%������y�-,��Í���쥪��@��8���m��;��
=v=(N��hE�}Fmu��a������g|�ct��N�@�-0�Qp�0�uS����E�����t��˭s�߶������v�>����CEZ��S�爍���WZ�{�٩�x�(����W�ߦ��-N��Z.�Ud?;j9����9ޚ:�ɰ`���N.FV��*�_�����2Ub.�Z7�C��e�	"Ur	�AX-�әa�PeS�_U(/Ԇ��LQ�M��c�	�wG N(
ow&{�NB5p�H�` $��c3���B�?�#����oO�
��RÜc�$�v�P��$��r��;3�+*N��D<oϻ\�(qĚ�AZI5�/��z�=�?W�r��0py��jv2�+w��k��s ���B�M��pkp�;ɍ����f�����.��(U���ZḦ́8������We����h",R��; ����!BH/����6)�K����T�$�d�u�%m�zH8������z�������С/�%,+�nV�bRc��Sj���y>�W�C��ے�vٺ�f�ŷ�=B� ��^����t��l�i�<Y��Y�
	����R����l
a�4L`�	R��6���7���&��e"p5������	_S�������MH����h+�L�]vA�E\ŠxLq��>^�n���y�KM<X_d������<%'�"D^]lK,�!�CR}nlv!4+��FV�K7Ψ~����JP��_�-��n��	��
�z_�S�a����)�V'�V�v��U~8�Y��e��::�M�a+���	�:�+�_�1������6:ϛ�H/(��8py[��*k�s&�C��Lb�[��IF�v��ݡ�Ǹ`t
2����� ����>��57}��Xv�����������.y��3~�z|؄�k�-�Hsl�%��î����ɍ�~C	�̜8[ ��n�~�*ؘ	��7IY�l��@������fV5���X8��RA�Z�3m��7 [�d��+���w	u��m~��%sj���X���P�X��|����[� �Pǜ���].���0y�jR.nn��b��I�����.�2 �$*i߃�����!;�O�8FdP>M{�~{F׳/��"_䘗qg{�P��]��I؞������d]g��j'�+�;�
�|�K����T���&U�=f}}���G��y͸Û��a�{nu���^DY�L���y�B���+Jk�NL.|�������]�u�
E�=��T@2��R�HjcR|z�b��6����Y��C�Z�Gs^�E�C6Q�����d��9G����R*u�}�.O}�?o���j��*W��ϠJ��[�*q�cd�U8��B��6 E�^��ֈGt��  `9�g��r�4�qV��R���
�\e$SZ�l�-~؋޲���^awt]ii�ޓv�z-��6#v�����R���r�y�C]���6�Vt�<ֹ�^��-���٠�T�SPl��t��c+3��%y��4��9����w���E�1d�Ƨ�d���Xo��a<K����jA�����8�R��e������s��S��)�����C�p�̚m�9j���޶@<���:���̠�\T3۟�#	�I��V3�[zf�K�B�/;T�ɵ�o�#p�J*$��t�(��%�!�t�S��˨jC&p��sfM���}��J�)���)A�Qy�A��k9�.;=�X%1\�y9��0�pPHk��j2��8u|լ��v�(KD���;[�m����rb��/^!d����g�[����>T̬�?��#Y�0��M9Z!���>V��s��`��h`��*F�(Cu��l��w����Q"h
l��
Tѱ'�C
Rg�v���9�� ��9�^"��,2�2�w���`�"��,�'ƈ��"�̹(����8���ٳ�FwX�V�G�K�jag4p�>���2O��]��*;dV;�r~�Rb���UA��1��~�J��B��$7?�F?X48r��H��y�F!����������[jR϶,�]d:Ь՟OI��Nf��L����D
�F7%�u0��_����?�U/�C<L���	��.��α]<��5�L*��M�+��d�P߉*��׃!��w�xu��HT�"�e=0����ļvƜ��/O�=�r?�־���4r�����9��#.��~�zߕ���{Hʈ1\NJX9�ȕ�&-���R��ݙ�*���,M|r?$l��I�-�����Ӕ��V��*Uv��U����;�$���m�NFb����<O�
��U�p��m_�J(�y�>���d��MB��?� �z� �W�$`������.2Z���j��zM��\%���B�2�]먜Uϼ�o�#��4���u���^t���o[ז۹.U�!VS@A�f(:,�3֙2a4v��d�W��U�\��h��n?*pj���ͅ��m3O����sϴ	6���Ԑ8҅"�S��2G��>@����x�1�`���髣��-ؗ�����z�P�Wr�C�`���a�@vh2<��9n�0ǽ�5o������"���ga���������aN���/�n���U�3Bj-���߉���-�<A���.;�@S<�H��3��#+1�5�3���E8l�"ȼ����	�Ӳ��
s��ؚ���ʈ��Ɠo��V�U�]������&3`�E��q�)�|	�hG��]	�'�C�o���s=rLCw����.�eV�~f ��d-,�,��=��ѱf~��Tq���D��ÿ/rk�Wo��y*�jO�J:�q�`�v4���m���� ���0v�K�4�8r S���d��;�4�M�%8����ק42��ǒ|�+4�XE�s�J$#f
�B��������� ��p�Q�֌{�5��I����}X���ϳ<Y�vk?��(��'��2t��(8�ڊ}�hԜ;�f�9�r VeLƹ�V�f��C�]Ә�B���My�WcQо�+dh�7�]�zam���X7*��Nd`���NR�0��}�#���Q�(�[ [SZ��i��-q� d	�KB�ٚz(U�࿤��㱇ߊ�@*(��5ء��+0qA�؋Ĩ�[�J�F�+b��:�jЖ`p�����V��N� G�pt�����5܏��	���R��c�6+�aV?Y	����T ~�G��j=�#�:���q���;�|ς{	�i���������q˓U�^%�_ ��ClT��­��˵��0���Qn�L"l���-�橅�A��>~��Sh�݀��z�1��﹌�D%���W��e�V^y|�9���s�/��˨_�inY��=�G�[���P�v���;�CsQ�dO���[y)����L�>�$O����z�4NJ�H����#���r��k#_*���E%?���y�K_����\�3N���U�/�&�	�`�2E��w���������dML�0������Q��
��՝��RW��/%6���$���b���)7��u�P*9U �QV
�ҼJ�1ry��sXlxV64EB    330c     9a0�����d*�e�E��9p)1��%\ҳ�yi�N5JL�EdA
hx��)A���Ly�i���ϙbj@st�N� �~� �� ;�F�+��O�0K�f��g��#n�x�n_֟�\-�
N�C-�xt
�x��c�i���{�иa���䨯�B%W�	K�-A�Msҙ��]l�h7�yC��r���/����&�Pw߷e���j�k���נ-δ~/j曟=]�ðWS��3Z�bQ����7]601Æ�{5HHJ,m��Z���J-=��:=(>��sz�'�i�w�^u�2<<u���x_�n��M+�4�(��ڌ��|�ݺ�z~-)G�8^�ie��q7s��N�&d+���6(�CA�w�y49�$ )QI�N���O��uP!0C˘t
E���Jj��i;f�j=��&�[��E;.��
����sB����<�D��:��|Ķ�Z'U�H5�Ѯ\�rf��Uc�[��ˆ�0�2�0����#�Jb謊��L�T|UoEs��w����jsy��}ءvy���B�|�ې�ϰ�
q�،4^g�5���� �Fu�_�Q���Fy2���&�"D!��8�^2�) ��/%�^��_�d�T�
'i��C��6�O;F��2��!�Qep���tX� 71W���)���w?��ްn�x�(�OA���H[¹�q:�.��O�8g��e��M9�>�H�z���}zr���)��\ݠ��*���T��C��]�V��=1P߇�B�0Ck � =!�������ǼG����tЭ�Ĝ�l`�p(M��m��m��Y�Xp�vu�e����1�j��k��<R�q�)W���{]	`c�M�IV��'v� i2 ڟ���x�#�e�l�z6NO*d�<��OVB�*�_����<�6w9J��X���!��eh� ��:?�>Ü
ߐ>������nb����ϮuF����D�>��:�����]�r��
������Z�0gW�_L'����<M����~�A���ϵ��7m�~щ��b�T)�r��`rTϛ�ҌG�Iڣ%M���Ȫ���^f0����)�I�k"�9��y"ѣ:�>=�H�g�P��~��3g�0΄�ma�8>��$4ͷ��,����w+��䯛��NF@st�U$!-v����/�]����Z��h��ߪФkҽ���S�����$�*7�����_12OG�A"�N���C��BO8����i��bz���|<9[3V|w.�t�-�|���&�>���JҤql�����.�.�$�ލeVw�����28v�q&H�p{K�=Ώ��mȡ���l�p�"��ڋ��a���C>��b�Am97pҎ_NF[̄�Q�e�㘐j��!�v :9�#��U�[B�K�Ga��{����5����WE�լ��oW4#�j��,��������q��+v%�s�|��p�L.���dj�zi3�m�/6P��r��X±.��|)<��.� ߶�d��4U��3��l��xz���$��\���)}Q=���q�+\�M�;�r���w��7}��(�')��!,�(	�5��j����\��ג.��=�m�2�$J�$�n{�'}����=<N+�CsѶ�lΝ���4^l��PѮw?p�M�'����RsRZpɶ�@ |E}qr��}1�)! �~	
EE�ӗ���f��H~���:R����a�fD�J�߳lƖC�rN�6P9[�dTѮˊ����	�GUw")�n����� �˜z��D!��LG w�T^'K��QKG�ţvc���;�[�� �dy�)Y��&��dY�`�Xم�hcA���{�h��Ssb܄�:=t.�1J+Kr���a�zή�mF�
���d=���
8���b}�8ӎ�`�	�q#)I �.+sj�7�?$��k]�ʓO��O�^�C3�Ze�	 �ۂrJ�pűM$诌���JPE>�w2ܰ�v��߾ͤ���HØo��_�9�v�RC�EN��r����=r�5E�uBM���/gZ�-�W����(�GT�ќi�c�)�H��?H�f�G�R� ��ƅ���06��c��fǻܴ����"ItM�-C��y��'/�$�?��\�^�z9��ɡ�~��s�c0� ��&,�7����F�G�
�1R�j���@g�W�zL_�"��Y�Tm�a��Ǖ���������5�I�X����b�g�VY�f�Py$����gf�C�A�xнz-p~��0at,W.����]�Yn��aW�7��������3t�`$��"rN%�1pL�:8~��09K����5�荌� LRJ�!m�
f��!@��Ҩ�2��n7)f�����~�K$b�8?�&� �}-��te�`�9r��"g˙���F�� �'��V�b�˛?f�7rP��������S����!��@�9�	McFWXRI����