XlxV64EB    15be     810������о�ji�,F�'�JB�ʦ85�bg�[���G����l��2'�ն���|a¬?�4����_�Mi-��N���PAkB��3�����,�l��í�SX�'�0�bT�~}\-�V������Gݖ��v�[�>B�� ;����:�V�?�掋�=�Nŋz"�c+n3#�J���2Q
S=����'ơ��TRH�ȿ�%m�����i��o�:�^87*ݕ�5��{�*؅�稨���{"�B�J�$���W��l�36��y��Ɔ�h��m;r�p�S=�[g��Z}C�L�T���#ud��}��9�Qs�Brm('g�'�~[��E�C3��"���X�5k����k���5�W�,z�)����� ���N>�/z�����£ h4�@�D`���-���e��ݓ;�(g�xAW�g�-q�g��Q�����_�9fesG<�Nx�ϲV��������-YZrX
jg����XbX|�3.�O8eC�X)Z��?�|�L[����ǭ��P�QÛ�o�k2!�:
�kZ�쾴kH����d�q�1����؁6{����yx���� �0��F4��w���x1 �+�x-y�	�+�]�ĵ�Vh�	Ek����v�+�"�x^�Ӝ���@��6&�M��f'�̊�C|�Z��BC� ݵ{����f{��YQ�0�dC��!�oc(v���8�zgCÛ���%�LC�2��!:����� ˠ���v�	NO8.I&J��R�ѪZ�`&�!�����B~����w�mV�4�f&�ɕr)G�޺#��J�x�S#eMM�K���t6d�x�.Q��$쾾��j���ϛ/w�b�CV��!�`"�5)����Ñ����G���F�oW<��'��[�i�4�y��ʣ$>��	�#�}���Mg;̎��Ed���M���e��+�ȕ�e+����,ܵ��"ԗ;�3Z��\g+��8�>�rA|���u�he�N�抮�u'�`���8m|�j?x��+�=ha�gJ2g�C�"��$k�ğ�d�y��qu_N�`�^+��I��7)���g�n|�7��7�Q4C���T�δDre������e;�!�$"�r$�u&U�l?p������C=���i{��ث��l�>/"�a��l�Ikx���(Ba��\7�V닎��Ƨ�jI��y2pi�=���3I��VP�&}���X}8���ױQ�`��0���Ou+�q����Ad�����CңL9[�M��0*h���Ѱ�l���w����T�4<k�#��s�������Ey����}���A����j��5Ff�3eA3b�`5�в�G���<�"�pA�x����4�z����d�u�UD2���ޱ��Ĉ'��VCB`j�T��i�t���H���9�~�h;5!i�N#����
�<�rV���TŜ�������0͡N��!!G{e@�q�5�YhDM�sCT�X���>g/L0�j��������r��>Gߍ�rZ�	��p�j4�P�����-9��n-
[��%� ��1�� �;be1�K�pBHZ0|˘:><t��7�����s	�"ʔ�OD-�M5A�6M���hz/O,��|�'��p��=}5z�X�>�b�m�G�tlc ��F:}�{����m�.y�P&%��O��T�Y	�,: ���������E(n�Ɗ�N���j�2�m%'-S��
گ"�z��  =�n	k�����c��Lw/a!I�*���nM�\�^V����੯�?�&���J)a/y/>�C��Y��C�;��~���3/�f1v�]ʛA���M��D���|���f�72O�
�X|�۠}�|.�׃��5֯Bv���sr�Ayo?U5����1r:���0G�SF�F���n�k�z*:v��d�~�N���'�t,�8Ig���M���u	s�����[�����$X��" 3��U�>1/�h	 �LZ�r������ٯ���e�͎������f�'� �s��>\Ϻ.�g����v5k�