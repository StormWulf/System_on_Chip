XlxV64EB    39cd     f10tOC�����'B��e�4ɾu�m��O����F�ʨ��с�|�����ѭi�C��V����o��-��n�x+a�Q��-��n��5�� (�SY���DRrty�6+��J}��DF4&���:�C�ޅE���n��v���&��EҺ�#ڥ�v&��?���B���.q�`�F�$O6{����D������X�j����.�38r�}��[�F�����{���~���Q�;UC�����W=�M;�$w?	�GN(z�d��#L�.�-9�1tr�'�=��mԗy�6�����3�O������3sx����lU��>�B���Y�Q(2u����y�b>��D=!���Yx״�PP�l����9�&���Bl�aEt��\�浽W�l���ğ�ycr��_�����pFq���^���JJΰ�rt���γ���^��_�}�f����Թ�RX�!���~�g쟬�d�L��}E�,_������յ��۞/D�E�lsb��#��š?��j�>�Q4��HB@]i���0�� +�g���8��Z�&��,�Ns���)��W�q����gv��S�m'�ߕaę���:,�M�jyps��|@�S��*)�� �q�1������� �Y}�1N�븏�+f���s���T,��{�va�B��`�0���H4P�OA�����ă����Y���;!ѡ�bxsZ�-���4� VG��Q��?��Ue�@&Fa�B�p���?w�����-��L%�Q�)F>q}�!�g�~�)b��n.�>������
A�_�8(_Tf�o�;�������d��ak�Y�Q��&wL��$�RF�6�Vk��YN��JAy��H۹��gm��8)�n΋�ag��F�r�d�
A)"+*E�+��W�`AU���kyh�Ґv����Y`4v"cT*����@�Dy���=ߋY�ʻ��~�#�-�)�}��;�JO�sڂW��A�����U�|w*�g&��"�d����g؊߫�Έg+T�� hw7n����T V^�\"�Լ�[R����bZy�1��T:�kU<`�9�+_��'�2�G��:}���c7�����al��q��ظ,1~ y�]����X�$�Y���ىG��S�N�� q��b��:.�U`�4yA�P��l�i��4��r|P9�gmۆ[�Vov.��:]��Y�x�sA��,΀d�='$ܶ�ʕ�[���U�>+hC{���	���ѵ�y髎��"�����h�[ۙ5νFg~`�UټuS
�����1��&�P�z�`e�Pb\؂�tx�e\���of  h���ٷ3��}��!=��"7nU��]��Ԡ�)�E_{,�*#�9Q���QJ߻���.V	�}p`����lB��&X��W�i�,��)^�R�N�q���!o���3T���1L�צ��hi?vf4a�C�k�����p��	�빻�+�ò��&Ծ��5~�Yr��L����U$��!��S��BJ;^�D�T����Yȡ9�,� � �#4r�o�m�ܚ2�(�{p@�+�����և6�*�$�ID����uAސ�$�����/��P�!��<24�I=��1I$J�Fb&|M�f$ՎR�@ۜbcY��*M
��fh t}|�͆��KCr:_1&%���1�D�3B߭�P��Ӂw�$6|7���E-�+Z%�ݻ�g(��oVL[�/�^���M8���&X�T �M/��}jm��́5u�OѪo���++��$y�'@���47�.(иf*Uf��8?d�d���JȬ\;5sD��t^�~��(u>:DmXP딱��$`�5�&M?��B�=����]|Rmׅ�7���ڵ/-%��|Ch��A�٥)�FG�h<��FB�wR;t�_��aD�&Vt��i���ZB{� �� r��Xo_n]:���oK���f�gf�4���*;�vO{(5���H�e\dB%��|�y�l�dQ]����.�4��AY7�;�k�"!�j�;k� )�ƨ
����L��_���JV�_vH����������O峠2���4;�7�:Z������ 87�<�h3z1�Ә���	1J����<x|�S�&��Oy�r��¬W*=*24A$����8�[�(O.�[��!Q�1���H,]��c��eA��X?�dqvW�δ��-E�z?<����>��&X�G�Dv������h�`ݥ�+���*h3�9�_ݥ䕩��Y_�U�v2��V/ME��zlT��r/�> ?��vww�}u����*cJK�����3�$��,���%A��
�����#��d��G�a^o�rR�if8���\]ބ-�!�ur�1V��+�W���S�o��ױ(h�i݊�Gꃤ�(+m:F�Z�-,��Ɗ��O"},�8��\��f�-�������A�Zi��e��L��h�Z�$�Y�>� ��E{�n\���S�b ��<?.qCx�su@~�"�0W�-�2��X����^T�;���<�7M�.�wd�"g�~�`nƓ�*�Z�u��hKw��ӀW�6Z��&�y�Foҿ�"��� ���=��y`��Qڞcb�
��S���~Z�py8� ������"�շ�����:���ҵIAԛg�Z���"JAs	{��l��#�X?-4e5!����$��Ԅ�e��O�q見�gR�E�̮����v�OK_b����<��ʠ�0@WJ����@Ӂ���"���>�Ym�����L���:e��f���v9�(����	�� ��������J�CJ�S�pIƽS��������� fhщn�x�
W��$�~���)5%����q1�&��j�rV�;m��O� �нyȱ�3m&T������Mqi��5�Ӫ�'5/���ݷt'�
`ߓL��.�3�
�0���#�怇k��E�y+��s��V��<�n�K�R_�����0�<��,�)Y�9\{k_�Z��dn�]�<{0p��?pi�{]"��x('�0��_�sm� >��M�̲GK/��I8Ҥ�4���<�׺���s�e�v���{�k��j��~tw�д���7
D�	��G/����w�Ϯ�!��)@W?~���xS�����j ݴ<�?�/��]� ^�!�
��G���ɀި��e��Iּo�SR}�]�>��RW���*�W�)aJ��+�*�S�˳���3��/H�ft\��a&���d���J���v��+/�I2%��������=�;�c(���Q��$'N��ʇ�h�[3_Pc$N{��%�u�YьP�e�����z���[l�}0�=� ���RVc��#�d a%CC�Z�i�m���t
!yI�K��E�;����i�Z6t�Za���C(a&���!�H��I�7WX-iT���	��vS�^��խ!��X�o�P��lM��^�be䙸�������sxɳ �e����h�O������z��8q��GF����6�H��M�\�0�$���Z���d�/K	��TsX�~�r�]�yd1��H[&&�~AS��&�񺇲�������P;�X�D�o �f���a�	F�X�\)�����-�P��m�,����̡$���޹�}�t
�6.�T������z�.Um,��cW�7��+I\���k��O����x'Ά���=�E�E���2>{9�jw���׺��q�h�t���D��ukJ��=0�Ƞ
?�L���x�G�x�;*�*���W|-�ߵlpm)��b����,�!�����N�ܯq�B����Q~�"����mt��