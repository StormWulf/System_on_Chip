XlxV64EB    244f     b40�3��9�� �����^<�� ��s�/�3$�"XV�]�^�<:��d��ǻ�D���`��ӡ�=Y$R�쟿!��^�2C��=�2�!\�����]��ۄ�N_q�l�6 ��=垇�A?O����r��`��U����;�c�H#э��"�J>����$p�0
5�k���� O_=�L��ۡ2]�8�S�eWڋ%���:Y�LM�ȘkܝB=P����ʕ)��V}:��ԵiN�l<B֙�s��Q�3k�� �_}�y����`�IPszr�w͞�� /���,v� IU��*o�+��u��)ӧ�ǰ�f'�J�~a�v��͘����=���vbl�9G����:�+��Y8Ĳ�,�,
z�N � ��m�.c�8[��������A��;Vն)a���N�y�/=�����k�~�f9�
�<k�}?�U�:@P�}|�*C�鱺���s^=�~�GX��IDG�)�d�(i�i�*G��[����=)J�9m�j��NZu�qZ�^������F�<GH�����Q����}p`�ǁʻ\�;�Uo�B!r�tq��҉,p�^?�(�x/�/����n�][�(
��T+.��iS�Qh�;��{� m=e�;+æ!�o��Ď���5�~�������k����e��\e�>1 ���T
���M��-L�����t��).�X?����8��͟�.	*Un^�`��z�H���	�D�8?j�9����js"��Q7`����-��@��,Q�&}��������ޡ��_����T����x�����z�ZqG��砄	��I�T���Hba
vL~+(����y��j)T.[�~F�u��dRt�S��P��K�<��m(.q��ZW�oY�'zؗ�^}�z,al���^�S��*3ǲ��s�G��BC�S�}�0fq�˩�)o;�u#�t�*n���w%�-mA��h詌�#���`��D-��{�� 1�R>j�"c��\�Ű8P�Bs��hL2WI&����^����O9S�e���C���<�:�;_��j�6uX���IT^�3�$�ଙ��X>��1��Rv�d����X%EԔ�"�֠om�m�-�dy>x
�ԅ�Ox�3������-�Z,CZ�p>�P��z�Q�p����D Й�&�ܠ��L:�4�w�w��
�P�7�(���6��u�g���R��5�*$�95�=��bh�+8����뺠}��F����A��[�7ܿ,�S]��Q"Pu�����Y����%�d)�w�M�b|!&h)�Lg�:�8ޱ�YXl���m�lC2�|k�d1��X�8��	�UQH0t�Kp򰝩�i��'���Gg�H<g���?P��E����vp�ۮsO���E��ԍ3Z�����pB��v��#�Pnmb8U�B�뮔��QV��A�,�g���_PzE��D�V�'P5e�X1�B�u?u*�l3V���}�H��'g��~: �S�=#IO���-z.X�&�̍4>��������-�!Xk���"_���犊�7��O�b���q�!�\��ދ;T�S����urf�JԢ����:��Jϡ���kZ���.�ƬT٤�t�N��]�b�K{�kJ!���9�TT{k3Rnb��P��&h�Pv�|�fW�Es�D�ߵd16��%<�#*Δ��hR�F���=��>
W���C�U�Cݛx��qN� W����#�ߴ5�)��]*4sm�#�n'�z|��q�,tgŁ��܃��$���:��wLoza�,}ܖg/���AH��$s�AJ���W6���Ǻqڝl]��X�g��.z�p�݀�w�;xi�(����>�8@�Lz�4ۧ����鏲�#��p� ��wG���0Bp���?1�frr�o��)�ܲoM}��Υ.�q�ؘ`>OV�k�q�C͖ͫ�ӝ���0�Ƞ J)K��>��ǅ���k���͇2:ns;�T9*�x,荘��`2r���tv����G{d�\�m������ì��������+$�}�G�<VD1��l b�'��2[v�g �����t�� �R�D���+^�\B����U�K<���۳�>>��&+��d_��$pH�n*�<W����/��XZ�+���9>*SI��1U���.�:���>�\�5��lv���#����X;O�hN��i,�3������z�y�%�[V���P�۲o����~�j������toX�?3H�
�~��f���s7p�B:p��A4�Pp�����;2͟�/���M,�Gd(�V�4� l���O)i��6�x�o�C�ӭ|;���'&����Q����]��CME[h4K��Al/a��&��㿪�a�j2%���w���0���g��i�˦'���GB�t�������7�!s75��s>_H�����*��j�ݣM�=��:��A2+����ʁ(�X���!q)!u:�"��	��ޜc
(ӆ����
,�4�&����Q���4�3� g����g����n�Ϲ�����8 y�T �'���%7����=���̒
w:���Gy�ǝ��>xs�T�~`�%q{ςwu�&�o���z=d��`-���;l-��9���\*/�y��#~R�}�ƾ^K�] Al�M73 F�7ȿx!��vȍT<H���]K����}&ҿ3���246to	�;n�T��9��6c�-܇�*{���oi�oϮ;�8t�kUI��\��itY:[W�f��D�����I+�[X����-5�������ᚳk�0��X��9̀�����R��m���r�}���9r�de���U|2|�W�B�2��/�2\��Y��