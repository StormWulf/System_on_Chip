XlxV64EB    1871     8d0d�5.o)&W)p6�
ٙ�&9 >����u����:�li	7���<:j�/��"G����U�y���+�����zh�Ҡ�r�H��o�A�3�+`Pύ��Q�P	+X����H=�vT�Z������މK�VpwW(�fU��R��"&0l�8Q�� \ ��{�Ts(�D�k��5��[/ZM�LRaV7ؔW�|���`nv��u~�O]������Ԫp46K�E��r@*0�"��VwƆ�����	5%�4��������_�σ���=��˗�߼�~+C��s��rID�^��љ�LM>�� i�m=��*�<k���{�Ҵ}��/��H��/e,�`�`�$�K�b�;qƝ�5���p�mp�ڱ�gj�)�ĭt>����S�.�- `�^�	[}��+���������_:�_��r��Gy]�ź�7IIɊ�!qW㳺���˦���K�z��[�>U�!���Ͽ�� ��Ī�5�絓�SRg���Ϥ�1P�^J#nV��`,֣Y�8����y���Ԝy_jif<c��H�T���Y���z�,�9���5	⠜VWD6.�IԀ��_�W<d-mj{�)�E�SP�a�dgp��{0��\��5U$'��0���xg(C?��*5�����J�gK5rqQZ�a�u������2�Oc��:���� V���8�+w�n;��~����-�_eX$�M!��3Z�*k�U:Ǐ�B��Ex���c$�A�~_UV�5�W�o����J�nۏ�0���UR���=U�N���!���������Ȫ<�S%����a^�z�[|Խ&R6]�E��7F0MIky[YFi���ELX����k��ܚ��~4^a^t~�`t�p%�����*w��P�5�6�z����{N2M&��$���5]y��H?�{F��ט�c:�+|~�����Ql�/�$/O���J�vJL�l�MF�ȫ�k��C_8��g�Q�>��@P�i�M�+�n�V�I���G����&����x���;�.���I��@.�M)�����!0P�Ч��3�K~����O�;�9	eʰa���
�`%��利*�sgc��?d�wKt����u�-
=�Zx��2�YE�+�S�auJ���7�&�܅hgB�a������Z���+	�d[tc`������*���V��f��B) �����V0�z�Ӣe@�o�C/��{R�
A��VX�s*~��KЃ̍m�z4��Tx�,*���iy�nGm5?bD�$��"�q��n�ia�X�|[�r�(�
�k�j�pf팳"kĤ|��i��/��0�5�	�(����C/�$� >N>�bb����׏�	�a5g���
��%,D�g˘�P�����@o�����
Y�̝��EE%.��W�B�{���cLM��9>\7u��7,���$�v��C�����G�Ax|9;��1��1�03����<&�Q�Vـp��u<��iv�}�)��b��+q����t&[�n92�h/p�A�_�<�k+
��W���}��IA���ލu�ӓ�<��,�1K:Iz��Yњ��� �N8�]?������l��K��5E�nZ�da"_���gj������ms���s!�C��U�����Ő���	<�����Y	vB�w�6@��R�}2���y)��s#M�����6:�h�G`ً	�n����|������ZN�{���g�V;�e )w`n!X���G�S�z�+�W,� *49�uI"����!	'�{h�5!hs'���-��^fp��\]Ʉc^�qC�	{���d����8����ʒ�϶��b��}��g��۔jI|r����z�\r�ֻ�=�(a�g�����C�%�.�������7�����\��?W�Vʖ���B�����k7�U�	�1��F����=!P
:�Ắ�t�k�鏪��|��o���oh��u�vB��Ijlht��$-Ĉ��Ŧ��ܒ�f_�oΟg'=e�����7�6��;�̙5xO�,4�x�Kx{�@�>�0����PZҷ)������y&0K~����<���(D09�f��h�JG񷫠T�=ҚՌ��Ğ"j�8Q��G��q�]F$�q�me�W'=���`/��Y��-H���𱼖r+˅[�!Q�y��E_���?��F}�E�L�N�t`��Z���;�R�W���t�>�K3��"bn�T