XlxV64EB    3f12     fd0���&�M�_~�b���V���A��Z.#�z+���v*��n��4-i�1le]���'b|�4QYWg�&ٿ���ղr<�@Aa�a���$�^n�%�4��8�����7(>k��[jB�u����l�xU��s
<,W�����[��%t��Yߋ��%u=�ِ/P<���.5Cs�lwXO��t�o9���*�u���h�x�Q�0Υ�U��7��G�gp��X�O�&d��*�FC�%"P�7�8��B%�A�l2��FqC*'��,=�POmV¿-��=\hl��������U)�L��ɾ�)H����a-@WU�f�j*	9�7z{F�����R�d��#�u_A�W��6�� &L���ً�(���w�Q$��v>P&�~���*6�W�`�ڌ�&7�3�G)��E�y�}`D!oQm�QӘ ��'�-�9,����u�pb�W�<��oQ(g�<C�Y_m�}L����Y���E�ǥu��n��(x.P����uXQD�������#����\�.+�_ ���|�lBz��`|xtk��J�d� ��X
���_�`�6
����'�������g_2>CSb�dFP�(Fs��
��E�](R� ��Q�ko�|]\ ���Q���'%9��/��̓�<��v�^���5�4���>�N NP��TgisW�����4��{�\�2���YA#���J������dQ�|� p�rāJ���a����ʿL�d�����pN���=�t�YsO�7'���`9�Q�g����w�2��=��C�,S,��&�X�X�(��9k��!�n�>l_"d���:�O�b g�t�D͛�Ǯx%�G�GSh��Qa|�,Vl�Z�?Φ�V���:䓦o�-d<���k%��+���#r��cL����7Gt[y��9FPF+W�+V��|�E7�|��>~/�����A<o�=Z�囟����Kc5b�����_#
��.���މǀ����$5��]U~�Si�0�s�C+�|JcR�.Y'����,�p�w�-&iFyd��=�P�x|�f4
��(��!;���94vZ�����+U4
K�:�h\�=�L��f$�Ow)Ԭ���k��Jd���sԎj�0�)7\�r��E�ƛ�'����C/��\�%Ba#�cFY�x�=Z��0EȆÂF >��~.����\��j������LwS�>�r7�C��/R*�}ʏ��[;�x?���X��.�S`�rm�?r�?��O�|�~^�#s�Ն�o-V�7��"�9� E�M�ߜ�7~JA��TPG����hm�ɶ~�&����R��,���4���Ŗ�`�9,��eǻ�fy��~��cē���sd�%��4^��H�|l��+4�(��g�����)5-:���L�P�9%sM�D����tѯ���g	2t8<��m�J�[9�n�����/��!K5������뮿�*@��yq&z��ܪ[i<�m>�_}2st]�(Q�;�o�n�$Aة��v���	H�Nip�Vw�i�i���bz���t9�"�xH	��f�;�I�V��ZĻf^S�Ugb�"�B�&c+7h*Xr��U;�lg���|]�`�����i�+��5?���"7��n暬��EAT�V��>{Jמ����	�GN�����2��UvgK0�D{G���L��M��8�Aq�C+���G�?1���q��1�Qf��OT�"vC
���W�2sŅ��}`�~�>�yt|�I��fD�����.B>~�b�����S9�%�DQ Ή�W8��v5�������˘�&� ����7�:5�#�� ��p�Xn���@���([:��KfU���/�)3"x[�V���)�*+��e��W���%����t���?�}X^ S�a]���$ؔZ� ��{����q��aȘ�(
0�2P�Y�ڱ���~�cs3���xV�=F�+KSq�g�@'J��@��e�����:\�0Z�f��]�]����3$)���)���5:*®>�[��*
ζ��t�TJ4�!�� �X��ijr��(#���1�R�y�ff�O`�Ta�ׇ�|  �#)�����6��08��ѿ����JWl\��k�3����S+/t�o��J�!�6���n���O�����w�{ur�`D����\
5]�8�^bD��j����Y��P��K�ӑ�vkO�O��'�W��0�-��g�U�"��	Q~V�M6i�9ӘQ��һ�	��fE�scx7Ѧt��-q��Z�/-����(E���^�8-����p@4�g��5��p�Ck��b��[�����z�;�k}ԩq�͉�>a���}�߆p� /Xui�l|@�x��xc3�H�4B������z��Y �o�+C��H{��/��"R�n]��E.H��7��d�r�DMȐa
7T���o�fr^;��]?��yd0$�>M��QgE��썄�|�����	�A�O3��?ܢ.�,��тd���'C�\۹�aYж"������6
����k¹�D��̕l�x��@�O��lݭ�5��K��q�#[,Д���	���`�=�phs΅V���}���ib���n���\�����c-|�*�z�FK�[�f�J[S�*Ñ��0��t> sB�@�)�hU�b��\:Ak0&��M�{U�!=i;�z�a���Rn��%��g
ty��,���r�����>:ϙ	�O��V�-�[v�d����L��Yǔ
,k��겙�{0�P4�)#��*h���#N�������+J��e���f��<R��7]�g���BK��t�E�]�lV�:c��VG�O��'�\�"닡xQ	L8����h1���S{�W��#_�c���_�^�kA֢�;3fc��Sy���꜈h3�,�{�%'��pĲ�U'�ˇ$0�IX���վ^�')lW�o�`*K!w1Ю�;*}}y-�2���+{%��a�@�R k�&���l��C���cw��RP��:R}L��QMF#7�v���Pe�0��Gb87۟��׹���`�	;1�^x2ڗsG,W�4)�s1������^a���H^���x�vC
�+�A+p��t�ъn�?���/y��,����k��k��z$tw�L8
1�5i�%����H���iqp�G�x�84P�,�|���9�ˑ�=�|�Y���{o&��HY���xz8�v���V��?�-)2�D��ER�@Z9l�^GCUsn�%�o�.?y�c�,�"z��k���߹�6E����	N�.���� ��$8SHc�J����� � PȰ6E��`�w����>6׬��'` ��,�bg Am�j7֌r�b�G��zօ���������|H��A���_7��6NO׍t��0�(F�ډ��ɾK8}�=��Cdd��F{	�/�����(��0�!����P��?2(��Tq�h��籚�S=(ʱ�V���k��,j��N��|����?,�ߔ��~XDJ��4܌U�x���I*��aT1uˈX�$D=�3r(�B^+��}�>c�U&y���W�T;/���]�(ȿ}t>ʼ��3,�f#�7%*g�x��n~D(�/��'�x;w.u^9���ip�?&����a�-���/�QG������Ѻ�,��#�l<����oŘv��m�*���IRx�쪸6���Iւߚ�LrQ�P�<��0r�b�C��&��Ս���|R1�ܭ��V�^[��a�B:m|���H�{ʕ�AT╝b��8M�`����YL��C�>�z󜽀�W&*�DG�$,=)�O���.6�3(~/�W����8焠���{�a%y�*\t�U�1B��3x���n�E�{���_�N��u�N����~�H�蚵�t^Y�at=�s���p�x��P�}�(�`S)����I�:s�4&Α�i��Y&u�G���S	�Sh>����@�s����s�uZd�^a�wF�0.��}6���L��ȬP��7����+%�!N�w2�W��|���N^���,��N�!