XlxV64EB    171d     860o���AJ�<��rםZF�K9�T���U}tp�S�ӄw0�:���*[k�j�2�
{����ZD����"$H����S�e��-w-ޖr�����Ё�	��B��N{��ܷ���O����	���0���%��2f0�����Vɏ?}G�'��f ��x��Ё.̺L��w���<nP��2�~�" oi�Sgb\�5���W9�j�!6�s��&�V�Q��³(J'J��8u��Hù`��OcH�I:�[���ϖM�_�ͽ�6ǹl�#G����6���s�/���F�����L�K��(��h$�C�~��u���7;�� r�r����N�y����5��ې�牘=�e�ᘱ'�D�'�������������2�%Ka�k2���*����sd���id=�"�Q��E�(��ڱ0}�:Ly�z��k**J�r���ˡ�:r���ح��4؁��S�H��$ ���X<t�z��,��O��8~<΁�6Pr��5?DK�����'���t��>Բh�	��Xi�vߑ{�5�����l{���ٓ�:�C2���ےl�?�$�[0Cj�0{�bqr��r���q B�"Y�|�H�j���T_aCN(�=�w;�j�j��3�ƾ�zэ �\5l ��@���{���T�(::�'��v]�:'��8?�K�� ��;W��D?e	�V�,��@L�����1�C�9ixѦ@�Ǵu��$���.`d��Q-8z���z�x[�I�n�z [R��G�e��@�F*����RD�������R���9}ۮ-�����T��T'�SxL�j���J���ɉ_6��00�n�狆�ձ2F ￓQ)I�O<�ϟ��^��F|v9h��f;rYq�e�AАD+eA�I��%���v��{Qs�����i��Z��Ҙ�tt�������~�]��9�q�J������Z�V�	l�)�KS�F���AT
��>z}K{��eeHy9���}��kS3.9o\��4���#U6E��X���P+ŕ�"�1LƟ��d�kv��k/���j��*Ѳ���)0��V�>	d�`�_O�Og���_��O���,�V�}�-��	�H`��oT�/�-i.�+F1\Yv�/=�z�=��?s&.a�|N�S�Gb���-�q�#�Ѐ�۱����a�d-'����N���ە���GT�F�bAL; i���|���[�E���%�X�́��A��0�g~���|���ZF�G8BG8�Z^�9���4+��"q���,g1��u�󓩶 -@)�w�Y�X "j�K�	4yp��� ����=��JPCE�hg�g6Re�ټ"�4�`�n�@q�W�	kn�E��*x��S�>v�9XV;�Y>��>g��%q������rNb���u�����4�F�*> V�_.�0}G+\���M6�R�0,x�O�S�xJB�vR�s.>���^i��7FZ+�9��mW����dF˻���J��ϧ}�\Y8��$��Ӓ��j��,����XQ0��]j�M"�|R3�1a��F~ ����7u\)�7��䊈���`� 8�����	d8�͆��Т\�����A��s|K��O��X���3��7"V�*D�[@\Z�䓯������k�Lt1�(�w���9�+����MIt&��p[a��%9N���*�M3���̚�x��s1}��-�����s��4N��7e��^d/hC�� ��	a�]jK[�*�c|2ˡ{�Ԯ	q���|斩,�G��+�J2H��f�)�"X���.�w4�#�9+�mF\��*sx=U�9��O�,�ɿ�
tr�?������&�ŝ_J�G}������E��G.-��u��J�e~����~��c�8���̅^9�K V�oCgk^S`�S��su�Fx$�LR�GO��ds.y���i�ښY!�,����{s�C�����<���9r���Fi������9�����Ԩ왡�������B�c}���>�a D)�|���Ҋ:.w-HC�%sE��}�:Ԕ"��ܲ�.V2w['n�gk�Z=�.��dי��*�L���3�ezpE��ɢ
������RcT�W�!���v�/��