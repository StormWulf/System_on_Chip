XlxV64EB    fa00    2e905��[L
�VZZL�d���:�n�q0>8\�(lf����~-�8���Q����M�S��2���s���� A�i���u2��})��>��l�1-�_�2�������X���;������b���k�A�LPT<"�v
��]�"��w����afg���I�L���I'�}����Lm��D���8��?V�޶��\�Y6��ku��|�S�f���6��C����()�^Uҝ�ZY���J�M��XUg}�ĶX�UeC'&[����Iؐ'�r��<����nGcw�0�����k�n��OЋ�Øz���Dg���1��Y0���풌���)6�����������%/A�q q�>�d,!9�e�m�^D�T�.90	ᢉlS���QXމ�9EZէ�<���w�W�����pļ�Y�$ƃ�a���Ǔ݅�-Y��/R�Q��p&�\��C��~)g���su�>s�s�b6���g�%Kڣlgov�4>��tW��7��Oʤ3f�ȿ�Tb�pf�1� z���עq�Ս���Պ��T������D��}�iNYwj/q_��eZ
Ø�uw�|n��[�ɝ>	?�����pM�.�ܬ3�~$5�b�����(=���ؓ�8S(���昂[�ݏ��+B�Cm��f��-J�._���y���$<��~����)-i��f<XE�WU+��3v�oc'���Z�▣,��%F��a��5w��a{�凯��zUy1��H�%�wi}Ks�����Lj���Y��
�j0m��X=��=6���ϻ����[�S�_�14�D����=��?e&�V1ܝc��:�,?�	9��T�kI�,A��~���\FY�j/�;nj�Eh�7�p�0�����U�d��e��Z�]��eѸ��W[ؐɛ�~��ɢo~�r�0���� �4����]�]
ʐh���u_e��SG�P
��
�>�!�	z�Gy��	��|ə���O7$6�*��*�+��E!�3U�.��h�jX�����>
 �-U��\3����<Q�&�J�m��#^`�8_<���b숛t�.��PȾe4Ʉ��=� z`�(�-;�_k��Z�X�$2	��Y�mf�����o��-Ka@d��*�mmz�=���}���ͬ�����I�3�m��^V�|U�(����
�;�T�P�"��I�De��:d5*:�j'��:��+H�o�]���K�mfS��\+��-�O*���"���Ӷ�1�^��M��^fv��b���-�*W��=YU�9to���r�d�4�i�w���.g�F�����u��g�ˑ�Tk�n�-��Ѹ��=A	�]�Y����w���kwA�x%�B�\mCK����d#���0���C{�r����vv�HZ@*�B|��̀����LJʼF�q��>�'��S�}a%&M\�Q��
3O�� 2��`;�&�����n׳����5�!~Nb+e��:1��~y�K�iZ�����U�3�(� {�$��>�T�������Yvf7��=k2�\vq�� <xݭ�N�;����*�x8Z^*&�w�����]d.��q��=�Ej��:@ޝ�kX=>��R�"e���x�Րx,[-�׎J+t?�O��l�����3	q���{�`��c����_�~P��JӝˑL��rB��^\�	k����U9��(�����F��1�Sp�:1�����䴪�o�S^'q��L�[")?#j�ԯ�D���d�AR�o�� �k�.Z�y�¼��D>h�[�d�]�`N�A�*�B>���,���Q�h���2���w0���z��?Ȇ�;I.�����p �H �<;���Wip�
��.t�7��x���ː��ADw?"��+�D��ul��ax��Mk%�E��1c�O���u��EQI_=�C{/dYW*� ���D`8���C	�]�c��qw�m�B<ⱐnM�x�$Z���E�#
@ji����z���8t����\�7G�݊�$�ЎTMxz�79Wd�A#v�����F 6�N_S0e�u�208E� ���cP�.�3)Bk�S"Y���ג�2#\�l7�L
��.nC)�Z�si+#�myq
xc��� o
�Q�m���8���ǚ�\�\����,�����;�(d�m|��3T^!��� ���Io�dN���,� ��L-8i^v6<�������oeX��B�}[u�$"3.���n�|bG�4�Q%���r��A,�� ���x����gp��|mk���N�k�Պ�_(�f��Cb�C"������k����H&G"��� S�������c0�l�G�_h�e<�^�d�j_����J]�q�b����Y#n��xP4Z��L���jo�O�$���DS�M���@�j���V��R��=x���Z�g�Q,Vk:�'�W'^�[S�RMK�����y��0D�^Uܴ�lz���}&P�:����@p�y�z�?���9��[�P?�n���ECx�7�av7~�-���*�CG�jH�<�S
��6N7�K�K���ſN�qԬN���F�
'ӻY�b���7��%b!L�ygh�,*��������*f���0i�5!_hj��|k߉��N�T�?x-`c��h�G����)����
�~��:T'����w��J?ػw[�K�:��A����I�"f�[,�](�e�Ɲ����G�t9\X���CD�qn�]j_3�O����G�N��#�8f(��:A�ē�D�w�:&��pcߩi� mb�tz1�v�F��)�E������JPrH�LL�a5�I��{�L������Xd�Z2��/�ס�F��Ԗ�-�R���|�X�H���>��+�6�6L��"/��Qp:���<�{�ğ	�W-���Upd�#)�ƈ��f��9W8���J�g����2
51�����S�f���ʀ�62��.�����ěOD�\�IE�i��XGV��"�Km���=��v�v8�X�btxOy8(�\>=yi�o��|s���0��<�V���a�^C�,t-t�g!p���_j@�6��v�$ũ=�R�S����%��t��V2gj�;�F�HY�Y�ۯ"�6]�ơuQX8��o�����<{�	ɦ���#�XQ�.���Ks��(p�%�m���J��Q3O}���R�=�_�������d�?�
�*�i��x�>�{0��&��+r�NZ��ɽ;�j�!��Eܷ��e�=od��S��sW��1�ɿ0*�*��4fb9�2����/� ��t�l�B�]�C$穔��L#��9�r2�Eڔ���0;d�:I��ZJ���BqL����f��[?Zn�o��Q"j�^�C��Y�����N�v��a�=����#�����r�J8��EX.�<}c�]^8B��ĸ�2�X�����ˀۭm��"�9����o���qދ����t�D9�oz��7�Q>��m����Z�I�6����n�Vd���wz���M���E���"��ru���B��EG*��p#2~d߳��,w���ÇQv�7�˞J4�d\z,% ���x&����ǉ{T Q��Q[r�ʃG�itZ��bc��CbX]��t��二��4�p���;�}5$�Q�(��I��Ӭ��H͗hm��6��|�ײWo�C�?��k��g�>9پ8�(��V�ˉ��~r�U� ,%Ǆq�������A�����{#��K�].����M����X�Te�o8���+b����)��%��Җ���u ��=W���2�qUְb>���B��:a���V%V�&�;`¦�/Ǣ�M��dC�$�C�5�J�Z��b���k?a���U�>����/�7꙽��EsK?��T��u�
�6�S<5�ʊ�u��e�~���a˺>��T�3�r�����Z �%�;�o6t��wU�f5}{�&gk�]�ZJ��N��o�Y���}��wh�E�C�+�J���3�ҁ���$"��%t���HVU�.'?[5����-�
�/��s�?䗇���J�ձ���L�b0s�uX�f��/��V�D�{�(��N�S9pTB=sRˉpsm��48�2|iUzӈ��:G������^��� '؍k�.1�ވ��c�'Z��+��͟ȔG�-����o,��L]�	��}���C_�7�%܊�L�^���[��htdA���Y��-e��J��O<��Y����d��ĺo�r�����{y �/��5B쳻���1���|6� �}ҹ �qn���m
AZ�~�p��U_����P�	e-X�q�BiF���Q�&r��1e��b�n���%�Bdl<U�V��C$�ُ�ϋ��SI�*0��O�X\��y�lP˩;��*��R+����s�ۨ�����|z�Ӝp.�bZ�u5�O����?��fA��e��՟�0bE���Ý`���>?nYU�KY�W ��(��-cM=(z��/���M�yyNx@��ꋬ��n�ç���H���=�����+���u����뤼!�Y"���k��~��kq�W�ӊ�f����[ٶ]$|��ױ�V��t�_Y�\�H;o���-vf�:w�@���R�����-u'�	��\�����P��
t.C$���Es/�S)�Y%����\90�ݑ��b0#����mW�]8
�Gf�`i������\l��9.�d�x|mڽj�[7d�8��1��|�5�b���A� ��PQ��{�WѶ�q@D�����F��|����BҸ������该���^�:�ݽnLPgu8=0Tg��koM>������D�Q��w�9�B�S��Q=4>_���Guli*{jͱ�Q�s:�8�*�q�n�L�݊#��ZSV!�1��mv���
�TE͸W���b�D�QFο�,�N��x|D�ꘪQ�#�ѧq��7�����B��VY�|q�
yg��ŸJ�AT��y
 �v���'�l #�3O'G��4�%��
��^Q�-{N;$F�~�)6��`�y�-o���5�b��®�&�`���G}�#mҕc�'���*�qsL+��i>`˼B�6�V$���l��e�sU��/���&6�P�3���>E$�s�\��L�'`���q���݆�K���z��F�1:Ւ��W�З�΢�?]�������������7�v�T7V(�G:l	=x�����٫u����z�@���庴�J,JY�����F�k�bi��S/�+g�P�a֊�6n�����@y%T!M�5��	9Ig�M;r�	�7N�@V��S���;���W�-C��,��>W��IH��.���ɶL�j�A���ik�����8Ν���Qa�)�P��aYV��T���;��� h��A,g���D�/�M$����6fg�Wϭ���!�\v�eJo 9MU�Z*ծ&Y3���L�HB?f��0a	B�Zr�֖T8L�E��w��x��طB��ݒ�	�]��'��	Ѥ��H��(�j�p��E"��Y���t7���ͱ�S-�n`�"���6 ��uo�0�OzL�{S�h"Z���	_��VU�](��:=߂s����~��Թ��А�40](^�oN2��R7�p1�]�x�P?�5��K��T[#S�̘�Aa��R:Zv*zgiY��Pe�+�.��_s�9 ��*MWb�p>=~bE�����$�EՊ��o�r��&��B�k�nd9��%��F1�'}�Y*2�7��qg��I���%g��3���ת��am�m�5H�Ͳ��~����aI6���5��q/��j2'�cP[�����2�kdO�J���%%r�0V�[7B���F�����Yާ+��?���n��Kn�ɱ¬�*�B�
cX`�X��3_5|��a��|G�d%����%�[�fnؠ���-o�"8T�,��	ZQ�����U��`���}�Q���S�i�z�oL-�: ��%�Ls������Ԕ S��kpԫ֎@I]��65��s�̷u��ƿR�Sy�|�I�~c7�w�R1��m�y����0� ��gdOg�����3W{�9���ه��ZB����e#��NЎ�4�p$%���vEU��=��� �3��l�]
pv�	R	E�C��wH����<��b�v#��a@J���?Kg"JU����Uq��#p��s�4�|���4`�wd׵�z�.B�Z��,�>F��4l��A�ѹk���Q"��/����%~r�����( ʽ��H�}�OtCH6K�wΆ�d1��,��g}NΘ���Ͽ�b	��YM-;�;��1��m���n�軭ɼ���A�&tͰ�;���'�@vm�w�CS���5_�
�y����t^	�5�Ge�Q���˪;>�ai'x$/��̨H3�g I��1Be~�MF{�k���(}��qU;f�Xc9yn�>wai��Σ+^�	�Xh{�$)V��v݅�]&�F��m��KJ���6�4s�$q�g�q�7X��]ga���m���DZJ�B�`�x�Ӏ����C�G1do��g�ŕ�/�c���mi�m�Ze��So7e�Œ���)��#�����My����*F���%}]���n�y,{*d��B����TF���	�Hz����k?�i���6�V��ʭh�wKr�6W2}�`J����=����W^p ?�����3>��f4z��,��zw<)p ��$�i񲲬N����`�A�7��7�Cj����4��5����U�j��kз�M��[F~�T_eDtO�cV�r�b&�TF��,���r��_��X� �rܯS��w�������F+n��{;�l���'AK;x5��,H�I����i:������j�!e�d5cI(E�3{Hr�މT2d/+_��V�Ŋ��X�(<� �iB|�Eǯ�dOi�X�8���;Ǣ�W�q>�~�����l�-��w9K��5��a{���Y�>0 Iko_�
_�����X�Y�۶Q�,?��!B4�L�֥9E�f���[ǉ2�T�Ф`��05������4�/�b�X�-&� ���z;4N-c�`��v��q�.�%�`��<�����+t�T�p,%H���䴎����u�'NГO�E,�;e� (���$�ȗZ���B\�5�,�����.�%+���r�AF}%
|�>��Р�꫺�@:�0�nG�$"^<�'�U��0���`P.l��-u���'�[�����>]:�$=�c:`�0(�H�8�B/���E� �{��Gu�Y�:Q��ҩj�@�ے�+l���;	�p	�-cZ=���h�-����B�4�G��gu�,��$����US(���d�ja�>}�TB�
�����_�L��8`
���I�l��`�g	y��|�a�
"Y��)��Z�K5T���yTϡ#�����!Ꮽ��5O����+�F�R�- .�&�xd%�`�U	+'��?X����2~�M�,��
N�Ԕ��F��� �J�i:�b��yH�Sw6�;�įN��,�#S����P�ǲ�ʟ���H��R�]\3�I��G�	��7����S#	���'V�9���f0ǥW�!��35X��q�NZ�N���Z����sr����ڽ�2�蘖�O|8��!RЉ���ȸN:�w]F��%]�H{6|��a�`�@2���9�J��.�;�3�!Y�~q�ŅE�9���hdhBȽ��A�:_ޓ�	��y�G,����~i�2��b��T���ә8_�w��b�Ț~�ڊ'Vo����$��t�?dZ�Z�̳��y�<]��ݰֱ�-Z�(`y�q����6�1L�Ͻ=���Q�NYO��ݤ��(!uo������e���?���J͜��Ԣ?�U.�oV^�"䔟���H� ���+Px��[Ø�1jG4t#_��NH�F���´��ڽY�ė����O�C�В�i-�793��F�ѿt���`�~�ʱ��v
*o�V.4� ~E�[oA�O�5- ��&��n��+��|��\O��ŶX��?h��ӫ�A|i� 0AK��������&��x�o!��=����6 grx�z.�z����@	����'
�Y�ޯ�P�>Jq�JK�9�ٯx��B>2t�24���>���ӡ�jo��Ai�x�ޣ%�yW��)�L�ObN��8%iګ\����
��;��zv��/S��xdw���976��d�o�/��>���QN��a�eD�FE7z�8�5g�"�p�MOŢȵ0���XD>	��m���{��jH��l���ns����#��[T ���;��`��u���O�^��>t�
y� o¹� iC��|�������Z� ����|AI	������Df[Q��l7#�=�}O�sFJ����m7��1����(|����|�_���� �n:���+"��[��m���$���s2�W|��9ず�ǵy6�2���8�L�eQ���yv1��wF)��H�B;fL*�+N-t����<�p	����Q�-H�P7���Ke�fԖrtL��4�j�L$_C���z��2G�ݳp��dOZ���G��X�1Y�]�q�i�ASR1�7���uk�﭅�ϿD��"��y$�.��E�.�j|;����ǿ@���i����E�i0�Hɵ��tg���#@�1�}��l."�7Vvc��]֜�fbw����F���ur��W�v������U���6��x-g%�5���H����jc��r�}ёQ6����o2��a|�����ɄС]��L{����0�/����s��u*ݖJ�ʄ�������"��0�/B�s�9��i�7�zP�X�PH[=X�jY����$'��' ��60^�Ҹ5lGS~�����|¨�tx)dm(�b�Ψo���z����[���|�Q�|<$Р���4��Fr�g��9<�%P>�Y�y�&7��un�W^_�f/͞��E4����%����C?������+׷��G�ϵ8Wt-m�)��:)&Ev����ܙ�G��p�����UtA6:��I�c��Hw�w��z'���k��V-����s3~g���;��|�_�xPj��h�'�{��Y�v�!@��ׁ���x�7����D��A�ͷ�W��9�kҦ���}X��B�㨇�@�O�"��蔛-��2`N[�
-6&�U�4&A	ڃ�2���T�8U�)w���].MS��>�ǗlI�BVT�x�v{�И&(F�K�Jg���ɨ~�����6��8���M+�O1��:�W��[x�&1e��@0K����ߓ����=�EHG�O��f�Ȗ#���ԆИ��P��F���͈��8��A-�9��;�]��k������>@n��
��V�C)7z��_-��U�~�^��[ZŎ��	���4u�C֎�vw�_8=N���L�i�$�T�E��]����\�o��J��J\v$�*)����D)��=�2�E���#������3(T1��G�:�M�E�{�~0��0��̘"ة5�#����RD#Bq��䡭����@���V����S���DY���4�HC�B
ۚ���b�kL��w �]$�P<��WCU�w�ٓ2��zt�o�M9�TOR��~X,�Ɔ�b3�>�j��?�t�.s���vE(dSa���F@�ګ���2~�ܸh9H�N��e��7�s7.��$�B5�������킋%��i�n�ܯc�_�P,s�u��c�k7U�a��߲�T@NW��6&�:�n��^�|o���J9�����,��I;<
B���+���vLj,�!3�a�5u�,��A^�0|"�g^*[�t/SPx���)�G"����A�TQՃ�H+�{ XN�E�!�q��1Wa�ˋb���J�C腆�S����*bUj�Gȭ��ã�Yw�y��
�R��r���'��dmMi�}���U����F���W���&Y8�
�`S�UK�%0	�i�i>��#��z��"��R#�9��^�X�a���[o��!Ɛau���s���م��}��x�Y���b���a�ju�L"j�Gv{��iF�e�U�>�񙅃4������fEm�U�$���Va�:���9'����0<nh` 	@�rAs'��byp��.L�.f�_!_j��zH�/V����(S(��	�['@�Ɍc(0b�{ȓ����.�_#���Y���֛��so�e(���J��7�J ��Շ��4�OE���Zu�:�F�;$���K6 �kt�v��C�A�J�c"���|�y�k�\�dYW�	َ]�k߬g�A����0�O�VUʨD�Qr	������u���R��ck�w	\nk�Ö��	<����A+�ϊEt$ϐZn�mE6����h��_UkR�u E,H�-�~��x��N�+��a&+]�^����� ]��V�P�&���b���qU~EF�}J���&��
<�dB��vEc�0]����^�I^g]MYT��ʈV�����}����_l���F�QG�)"�s�o�!�e<O�X��W�8ᕏa�dm]����I>ݧ&[\M�]������Ho�d*5n�	)V��[ �l=r4��	��ތ��/E��x����ga�N��Z�3ƙ`��mf�(����w�5NHА���Um$�#�P~��O�i]���'�G�;#<�3|A����H�hq�}�Z�9�������q�=aU!W�{��Q�:��p��c<�� [PZs5��|����-;�����˱.��^Z�g���x��.�� i��<z�����Ϥ�x�'� ��=��ڃ� ϐ���?T|�����$J��EQC�s��L4ɽ�ט�iY��B._��6��]K?�E�[j9�r���N��/⿒Z�ֺ��f��CG~��znX�(�͆s���W�K�Ï2���뼴���!\=փ�3��,�5��m������L��P�|O|�qk3A:m?{쩆*�$�] ٨~��ɼ�7�;�zNl��~��QjC���Ij�uylǯ1�N]�2yt��T�<�뎂&��
�9%C�,O�V���^l�� ?�ؒz��g�������$�;�o�z������jE��9@�lq`=�M'ru��2�����%�?�M$����3}���İ����rG�/��`x��Q�rÔՏ�������� CX�5��#H"�897T	�{�l���/� ���X)�����yح���v>�X*�h�F��Q����pP�|(��&�FɋJQ�g�L[ڍN%"�e�UfR��[K+�m�d�,Ĺq��G�?,��H�lg�a�q��ŕ�8ӗ�1L�9lNz�n��aj��5A�`�h�o��ˁ��)��k�V�Oa�/dc���s A��p�}DdV�Sݽ[k�P�عPvL��~�7��'^�?
���0HS�s��F�� cÂ���f=�q�ܬ.V\1X�8���皡E���ڨ��9�d�{��B#h��؆Ƭ�V{�	-�m�I����h_TN�;, al���ta͍�Ï�{;��+�7t�Yz�=Dk`X�L���6��)�mj����R��y�@xYa�Q�We�-A�-[���T���2���1�p�P�����۹����2o��*����]�� C~~"���1�T6�c%�q���A�R��t1�fi�l��|���������v8 �k��D�����_v�e�X0��p%����ɓ�f��В��Q�>�Ƭp(�*\V��~Iy�B�g�Uk0جy����*�GO��k�������J&RXlxV64EB    fa00    2bb0�;^18=�+.��uH��@��q`N=G^{�a���XQ���:���\�)˹F�$To��Xg��AgP����¯��a�k^��F�I ģ	m/��1{�-��.ѓ�1�����r���C���xu�)�V�����֊�����[�N�>�,���ȏ��W��7*�'��eU��w1к<�VQ��<�>���ێ7}���8�u���=}�1�\�>c�v#6$��N�.�vV+с[��b�@����K b'Y$��_ޒ���,@�pN?�ڴ� ,��(I
��d����۹؅6~��ߎ���G~�K�<ǛN�������;��
~qnBw����W&k`$�D}�bb���35�-��E��>�e�`"�R�*hܰ��G0���Kh��sX��TBmG�X%J���fio�ղ ���4�Z5�j�+�A.#Q^�y��>��5�󇚦�o�F���?�w����,����h�MXg�=�a�
�t�(X����]�T|�Fu���m��%oת�?؍�skc�.P+	�a�z��{(�3�`Rx�Za��?.�i��q��]�K����}����i���$���v"z����Ul�Ә��`6�^Zy�W6Z������>�Tj��_����T�/[k~Y~��F5�kC&��m&۷�~�ƪ��ͷ�R*cC �z�~�z�rz�	�R����G���˼�z�RT`�oҶyt�˥�K��޳tx�d�ub8V�"2�f����瞆���_�d��6��{ĔrgV�ߝ!Qv��q�M��q��.�Y8��`�͍h4�����)��B���f:y���E�X�����˼>��k�=lvޠо��#Cq��`�_7�%��������M�q�8�|�5�e����%_��]�U�\j�7�+R�����n2�������im�I���A���ro}�*t,���v���jh��R��M���4����Wu���T�����=�<	MF[W�:� 4Ŕ�L�g��/���Ͳf�$ה2ۨ҈�~����T�>L:ܣ�R�@��*�X�eoﴞx:��n�w��=~,���Pzf�u'Gҥ���Z�)dPh��3�x��h�ъf1��ej~�3	�`�Ę��
�@辱�?����l��� �����k�Z�$�EX����v{�I"�����-��9�kxH��ʤ�Ҳ�ޭ>K��:^y��;dW���^>k����!y
N魻i1�[�;������j�1eQngI�bx�`� Y�=��DB�c�qKג�M�'��G�Lz�Mڽݮm�?�	��4���3�*iu�'�������"K�ύ��ەyX��v���Ms��h��lY���x��E�dT���8�' h�.�jTZÿGM�V�"�ĸ�a�=�n~�%����J���q#YA�bvԖ����:8��80���d��R��~����r�L��39�b��m��1�t�O��.�|b�#h(@�s�=���'�������Q�A؎i�I/�*f`8G�`���iA����m&��A���e��8h����f_��>'A��'#θ�<f�'6ޕ�94�;�M�Vɥ�kf���O:���?��W��n��O �F#��V"�ʰ�K	�o#���`�􋒬�nY��a�E��}�y�
6���c.�"�I+���4�[���dK�Ŋzz�f�$x+�i�혔��<���J	F��<��R��/�������2�#p@L>+�����h�M�VSQ}����ڦ������K�T�P��%?9��?+��%�,&�Q� Oҋ�RQˑG]�5!�aHt���ȃH dT�0�,�CE�m��fh�͢BK����c��R�$g/���X��*�'F�p��A*s�D���W��]db��������_�_6^�)��N� #��O�[uj�~�}X�\ę.6Q�/�����-�k�:MC�����h>�*�1��V�~u0�ڭ���W\�q�Z=��PZ��?!k�-ݹ��)�5�
�*��������������ۤ��焑Wr�#�E��Q����ϕ���d�I;�ʕf{!�9�Z�u�	�8�CQox��=+�tP���@�#5���Đ�v`\k`�!��]�D���Rhky(�����W̜�j�\�Rno\��z\jĝ.�h�]����C��CFp��z}�� ���؈q�Z���Ŵ=Z{�/J��N�I����	���_��|�M'�c98�c�;������Φ�L���Z���1�n#�ލ���8�$�W��J���4�Q��F�}RĞ�����KP#ĢIN���3�M���n�)N�]�v12�����P�O��s׹�E�&�N�oh��&�j$�0Ƨ�RN���^(>�� Ds�|�?^�r�}�Kv#��k�Ƶ��r[�3a���Y�.zw�b(%�
+�H�孲/��g�\-���kf'��{)��FX�ic�`=�/J�u��
>)���~U{[�Z���UA�+<��IG
ܝ�Jh�2,���{*&d�2�D��f�P�o�)Z.I�4�u-�/�Bݣ��#!b^]6��GVQ�$3�;��#���_����RL��ֿ�2�
/&u�������0<��^��	 q�X��{'*9��2�r�oX���i�T�2h���vj0A�:+G����
��Z+�-m0G��`���#u?���w��NxRh�G��͔T�t��+�[�(X�t)&�#����)p=�!��w&9��1@�͝�3�Φg�U���4�K ǼO.��wi��� ͐��J�x �qWa�r�A!����p�X�pC���w,�rDs8�^�4�pF��X��H�>a�r�H��Z[qFt���o��%�^���n� ѣF*<�vN}�����kz����30���W�#�{Ȟ>����� �����gh쳳��d�g�8e��=d���	\Y�G��;	�%��H ���;�M�DjL��l0D�Ɔ�F`_�q;�1wP8=C��Y�r��'[?��	� h�V'b���ayq�X��$�LLA�0�=�HY���[�����]'���>i����: �~�\z�B&FU^�7q��:{]&/�����N��|�Q���*X�VH��)c�O/���?��ے�[0�(Փ������i�R���ė9j(�*�i�P�;#(h����{(�_��-��6w���&3�:U6		'�I(C�����z�fM���u�A��k0���J���ڤ'B
I��Vٙ�:pv��{�@�EI𙱄�6	�vF�$���̡2掵���޵��&X�>�:.������ɠ/x�x"@�e*@��xl	U�9�u~Lp𷣦�m�h�0�ǩ��?���D�b���gW7'��e�o(
̏�ܒC������\���ҫ��V��1Q���I�3ZEsR'�EQ��M6�|Qɓ��ǔ�5\ҭ (�������$�L���D.p����$e��PI�S�r�"YW��Z$�[N��^ˬV5�6h����W����� ����̕ʥ���/H^%��U+"�E_J�j�����Ԇ�;���!�e�k��z�V��Ib����Қ�z��6=���N*��J=u,c~��Y�e���/B���`�b�	��^JO�^�Э���U�x�_�
q׿��i_ -�b��i�$��?B�s �̓�[���W���
��~iUw��G�t�)�zkV���>�%�b��Č�S�)���Rn�d�s���+Ǡ)ԝ�l5��Y.�M�ϬB��hY��6��n����iZw�'�],s �Bm@Ix��0��&��axX�/K3X55-,pj�}�ο�X|�&�$�[֩��9�]r(CAK]q��0^�ly*L.$G��ߌ����=�T,ȇ*Z7%���hg�!4X/�_귩v8�20傇H.����IE N�\�#�q��������k��� ћ��vL�9S}z��&�zF���ob��yT�./D����	sr��؏�Gސ%�V7J�@���§Gy��Y�L�W�l�RB�,�c����mnOtϮ���J�ؠ��Y��*V)����G�U`�U���<�<NJ?�j	�^u{>�����y�vZ�ʹ����u	��邯���"�;��[+��Nն�{�>z�ͷ�`�Ñ��;�st/t���D���UΗ�<H�?���� ��br�G~�m!�y@Aw_y꒤���Vl� `"3�9�̤>�҃�bn9��<��}����&<>x�:�)�:��މ�#5�?89�0�VC��ǳ��%�祈������l9j��4t� �}8��}�,��*�π����*��rU޴���3����3���s~�(σw�ռRS���̅Vo�����\L}���2�_�O!�����dß�_~�m�U9}�=5bXI��S3�Q�����UyjVyy����tt)�����b��3���_e�b�Ia��$/�j��'��4F�2�#ň�����]0��C���+9f��~�E4�I��/aΛ)�`��V@lb����1�יD�7v�	�z�EH�t�EeUD��\�u��4�HV�q
)H��;�I���Q4J	%n��mD2����{;�%'����J�
�N� VO�l����x��50͆�)xdb�t���]��@-�i�p�ئ����d�~$����^�������TAg<��R�1H��l�s$��R���V���`6�v]�I�b�]�R�K�O�ŀ�T������긛P
K{d��~�^��LNS?^t�M�9�v�u�j�� ������7L��sx�W�>��0c�c$�/�C��y�P��k�C ?e��1��P�mG6�.�i���wj�v��K%�����$G�k9�8�&W14���0�`��7�a�w����cM�Ig0����m\u�$�lݷ�M/�!���fP��ĩ�m��Z'A��߇n����m����At3�	���Qh-T$�:@U���⠤El���gM���M�����~	���a�6Uk�K��~��b���ۧ˕����]��"B�![�%7𓮙�$0[���H�tL�}S�jv-�{Nh�0�Dv���]QOJ���K��&�%�,�u��dD�/�.���^p2D�m} ����L��>Rar0=#l�g��K#m�E�( _q���,�wI�Ng�|ط�+�mS�#-�#~A{p-�ѹ�z�%���Q�M&W����e��~�~L|�Z]�P����̼�D5����^������ȏ��w6��<���R�v>�t.�<�[��a�ZJ�ꩡ�(�-����`���3�*:g^�x�=v&o��@%xՉH�U��ʜɵ�VV�Ҏ�����1jN'�s�7�>�J���!ȡ3}T�YA����F��.�W�k�t�h��A�yf�ߕ�Hmv�h�F�P,0`X���u��uؔ�L�h�J�X��x�/�Ǆ��_���zQ%�]l�m�o�������7����,S(��O�@9�(���C�s#��(�CU�Jb�6t��DD������k�=�Յ��O��a�:Mc�m� �~�K�H� �>Os�#���_p+���gN��fQ���\��֍W�<:4}���j�}ul�7��n�Ѯ`�S��3�%��_����U��&͐�y����P"�8��*��LA�˅*!�`���x�}�E��Fq�6�T݂qX���Q�����mTZ׺�L�)lH���8�C�<�ȷݙ�((����k�>��i1�{����RH�͎���6o�Xq@�g��~�j.��{N��M�D�u{������`�nc��N��]H���o�/w7_/qI0
'��]��/��_�����\W{�Zf��~�jW)�:�k8��jk$_ʜ)��R�&�<�L�\�]���1�T�^�ǫ�S=��G�������!1��XУ���z�W��@1�����1�
G��`�C�g�h���{�;��ʢO	5��Գ��"-�A�� b����}L(Xk���+�@�$�,�|d䅰��aNЀ�y�s���uq���2E����+�%��@�/�k���bs5�_K��=�����ĜU9��D)��7ϳqk7x"db��ᢇ����8
{Ir�jq�Ҏ1���'.�k?pe&�稲�B��=���k�lK�H�p<g�v�2�,��z���Uuav�.Is���ߠ1���*�P��ܢ�f��9��B�n��ɩј����łH�1�촥T`!��@]���U�� ����at�D���!s\DA͇C	����M5�
Sb~�K��|)�)�i�C|_b����6�
���vFa�	��?�|>�,sˍ~�R-����vJ5�{��W2��@ӱ��@v�GZD�Z���=����z�Ip%�$�*��첽+�n�������n,
�U���}���A_�*I>ϊ~���眧{P<�������jy���P����u�aպ�� w���;��+�䲽�q��<�#���g��w��L�:�3���Rnj�3�t5(n%��ʥ�����ɓ��2|�R8���t`&��8�x�x&���� c���u?͜I�!����mS-��OP���v^�� S��m̷�-e�*8�=���u�ܿ4Z�\���)8�=cl��d�=ZI�˥Hz�� 1/@4��ђSF��+P��Ʈne�~���v�^r�L�F�=1���d��h�I�'�����Vc�ݤ�đ�y��睖��֝��;ǅ�;Z�.5c�wɎ�������y�1̛����,H���g���g�֑a�O�;�|a��Y�ނ{���{ ����hzVUR�~]�
�7��L=���F�nƮ0�yw��呋���#� !�������y5�݆�L�}��Oj�����xO\K�Ψ�~i5}���Wk�cǳ:���Bo�*jQ�+ʸ�����<��l��.�)�Y�Z���{���Df�4Q����%��J��VJ����Jw���ߎM0mĩ����OQҫsE:?J���
��;+i�Y��O
O�B�����3���6�8�b� b�!}�n*��>�F�	z:t��V���w
�+���j��q�/��f�}w��u)�tN�Օ˒�o���0�
lvL��9#��0�����a�%*�oo�|��ӌ�W��{��$�j�J�䇛�g��������˗��J��`1b�7M�{���_��"��m���8�x%���$!���wQ�!,i��DeA������z�N�Bo�Q����/��l��w/T�L:����-�|�T����RbO����U�'k=���a�Ш	��.H�a_�ì@��荧�ʯ�>�#�iV���zN #8��u��nEK猴��� sp�֨]4	PĠs�%�y8%x���v!ԟ���w�� $�r/q0!D���cGW��.l�?z�=G�h�;I�����č�+��[w�갸4��0y��L���]�6�b1��N�;?�e�nAhsi<��9���f;j���@��l=���Z�s���v�>�ib�	K�W��{�8<H�OYN��
6����6�h^���� $���G��~&LG��S�=K&��$5}<]P(��V���7yv���Wx���]j�6۠kZ;i!Kv2��L�XG�����W���_.�\��
�9R�5��|?����%�(5�b�����[�,����������/E� ���{2z�s;Q��\���Q��u��:���bE�1\�=K��D;`x�Ͱbs��9l��a1;G¾���*,@��ؠ8�=W~���*�e8�G�Ӣ�W[�g�b��]�;4Y�b\�XV����e�4��Px%����'$6�ߖ��KS������D:�<e��(B��T�t�B���{e��+`Cl�^���
� �G�x�������}캩(�/̗v2�( �C�hp8�SHw�Ix3�ef�+>#���N7�\���c8���e׺ܠ�9JUO���ɝoI��� �t9��6�4Qa^*��5�W5:A'gJƶ�x�N&��}�o
���v|xŸM��T�F:3�����!$�G�������\��$�}n��'� �]B�)�3�S��� 0�Li�= �>j��� �2OI�iA�&��[��Q�s�dKKFFXβ��tO{�X_
�L��hĦ,xW>� � ��w�2�T�q���RZ�dH���y�"Jb�����3��Ĥ���_*��?#�������E�-�j����
z�(�#�����#�7k��"�V���0�ad6>�1Z�?�k�hcʞ �g!��P�SH_/�$�����f�ٮ�j8��hDl�rY�1/'rj�N�Wf�a���X��|��<2K�@��F��$n��3�n�����=\�]�f ��������MUBw�Y��)� ��G�q؂[	@B�k�R3�mհ�os(�ј�թ*�X~.���V|�Ue�k�iwK��}���ђ|�)�sif?1����	�-0WQC�5:nb��1*�	�����Շ�ω-�,vB%�$�י��qf̦�$�)��[)�>��Y�2n����'����9x��r�R��^G�s�pq�~��ē�es�_J��gVv�x?���'~��j ���|*;���뙜��cHN��?Z�O��Z��
C*u�?_��`B7��.q+��(x��EPVH���nL�9僒���)����KF���I���ß�A��E�pi|"�>�D�r�ݭ�X6��Nw���31]Sd�H��i�ڣ�O��˄et� F<��Њ��Po7�AO-t��B��ZΥ�v���u�K�3��8J^�lJ��'y6E�-��U����͔�N(s�w���b)�Y995��S_�I��&�a����ĚP�}k
�%ǐ��.�}P�;���~Q�]r��Y`7�x�vG�M�H�����te�oLXE��:r��҆?�N�@�q~�/�t낙M�����c����ʫ
�o\f�VYy�z�����f��-!۲O´��J��-�QN�a_�`�/t�ڀ���i����xZ��a2ɋ�#[�`�ע:R!FBQ�&�9�+�$�Pz�s��j���saPQ�������j,�\O%9����U��etv�CQ�.'�(��$4��y��q'[�����*0	�ƛV�w~��.������ ۴ճ}��?������I��U�r%>DH{%B��<�L�~jPI9�T3ޕ�CsuX��`z����и|,Z��j��X���;aFl�5��8:�����ߞ�Q��y�<ђ;��"Z�$�>I�3<�:Z��� �A#.$cL��>��gU����ݺ�i�T�ł�A� ���U�$��9�LB������H����ΪZ�<���pȠ���H�����h-�{� �kD�j����/����S��WBHoS����C��3w���'�Qm��z��g�T���s���у��ә|�z�XH*��	���3��j��w4Y�t֨y�3Y<�WX,�T.e�9�֛WZ.+k����r�p��P7䛖�6�\��X̮�U�ӵ]^#�s�-�4����Y�a����]�Y}ύA<�&���7%���<.Tl?���i2�)�/3!���8�5����-6Wp6,�m��ͤ�q�	Xa\ETG(3J���h�Q���}�3��C����%��t�~����UKM�Ӟ�-0����s(/F�2m�\�����:�m-*�_}��ӝM0	��YJ��r��G���Z�\�f�Eƚ�m���`�?���1c�u�t�Q���Yf�j�Î�J��7��c�w�:8��X�0*T�YoA'�t.B���1��X^R3�sg�G\�q�-�k`�n]���I�,�>�F�����l�M�c葕%��##긯Rz�5�2o#�x8��6��@�R-�¡���ι��G/�>���G_�o~�Ǝ�Kֽ/L^A��%���7��N
S����ݺ��5����9�>縊�^>�o.��5�����^���8�D�p1�U=�cӠs~�" �������E1�\��+˓����ޛ�ֈ���z�r���Ewy���At��� ��$�wt�X?�{W������\- 0P�RH���� ��A�.�x�A&�``���@�r��5�n�h��v���3N�D��<�d7����9�t������[��#��Z�����2�;�N>�����D�f\F�!�����1��, `�y6R�.?�p֐8�qR� ��喦:?��6�H�5c�F�6~wc�,�!���Ɂ��~v�R���'xW�i�$#B0��'��$s��j�"Ge��ש��u�k�_oj;G@䪀T-��2kG��g��@<;�h)odݣ󎶲���>x�1��%�}���H�4V�7p���5�bTy< y��p�����MA6�.�P����ɬ�'<����a5�3��N��%���|ԏ��IV9�FM xP���u���璫:�����ɳtF~
t�W��MK����xd��dwv�1HP�+�8�?筋��EV[m�-Re+�MD~4��"��Z��dR���:��~.\��X.�a��e�mIU� � ��*56�� ����ɴa���a�i��'n���A@ �'�Uh���ʚK
J��>_,�*<0�Q�����ס�ld�r'�(\��/^�)��8i��ӧ�����߲m���7�ME�Wҡ��h
�Ct-V��hC}�'=��7m��C��{N֦������W�k4���>��J��9�pWSl��s!O��v�� �Q�`��#8Y��3%�K8h���e�B��G+`:�o������t����
e��Ч��|��ƃH�d/�2͐T��I+̳�ncp��Y�����Vъ)��i�f�S���"���{oF!��Tg����rO",����呙�>a�>�b���D�C!����)z�&gk�4gC�/q��IH�et.P��V���.G�YIr�݈�t���
7d� �(����c��C�b^9/�<+�/����FZ_�g%�7�*��̝<]	XlxV64EB    a433    1bc0E�M^ʴlg#�G��,����L�se�xM��rԠ��"wj6�D<d�p�c��{��Y�D�-syd(MOvW���UL��-jY���֯��q�u���]°/3�h1�ۥ��� *y�9�f$�����v@T�K�e)�W����`%�_a�p�2Gd^CB�~����M8��.z�����F5uNL�HJ>�=�o��"�s3���ئd�5�8r���pK�ܰ�4����@ӽb;���k��q3�S��;�O&��8�K8�q�:�r�ej������������T�L0֭)�P����
�J�z���hkLu^����6k�� ��.�����V9	�/lrH�Y����Q�<�Wߌs��)�/�_���l:>dVP�%��i*RY��&>�%�� �_��Jn�$�=�(�*���M�Q'ӧ�s�뢕�N���t�riǓ+�1d�DC����v���Pn���cP}� R�!�v�����j��L,�������>�)���8� ��\�_�>����/t'�S�bصss�^
�x���t��0�8`��n�To��!�רX�j��)�JWQ,�&�Cӵ���ފ~`q¡_� KI
3z*^tC��X���FM&O6É�n���^���-�F�hn���`Ĭ"cE��x`�ơXSr��ONQ�1˗���4�w��놿��z�^)4Ye��*��y��Q�G7t�U�he��B�6s9&�4Y��K��-A���h)���I�./V��Z`���e�����z�b�o,�u��4&����p���p�+||q�s�PD�������a��qLtT1�h��$/�g��\K	\�iu[��q��ӲJ,�%�ɭ��{_�@�:h���Z��Å� ���Ù/����|b��N1��g��n��de*ɢ��.A���9 <hvҧ ��/L�'�f;�����Ʈ�v��r�qC�����e0������Lr���%?����u%�"�����&*�����1י@	�l1��k�����k9õCvy�˒���xBG��)� �؈�H����x˳��~�ƀ�D�~��H0l�w.�5ĺ�0��C��򤊠oչ�h��B;Ռ������?�^�r��6�38��x��	U~�6ڞD5��#��& �����׍v�֎ZB�h��4 �*(-9�$�˫ ������T0��b��5�� 8�ߝ�SR�^B�(O�,��ӫC0mf6�~]�q;���b�����u��1va�����5���A�í�c���v�)B����[t%F��&����<Ԛ���	��b�r��nٿ搔��g�E�Pz����B~M<�@���b8�J��RZ"�z��4�jɢ���
~*�p��xD�r�����ַSq�����b�3�E<�����o��f����C��rC�:���3c�؃XE۝�Ǉj�݆/����R��(pqH��1���m�J���`F�cnԇ���5�)��[�N�{J;���� 6�_O�q�5mɹz����ԇ5��.֨����eoD�
��XGd��?�q_�n}I�n��P�G�|�W앰��B�MԅA��9v���s��n�h]�l���_�� ؄.N�]�>'�g]Q۹�(�WM�:��?���˳��r�ce�[���oK�&jE�-(_��.|nRU�X�|-���E�w�А ��;H!�ym��N�+�w��>���~�)��u�uZ�H�����tUd��
���u�l3,���Y{ �v��5j�e�˘
�(`�n�9�H虇�� {�Y�h�TS�"����F����!���vz�������D`A�n���yE��-}`EV���/���ԃ��DU�u?�i���,J���|�p�~`�>i��"Q|�`�����F��x	�M�ݗ���g�2���B���w&$�� U���I�����&�WrK?� �4gX�/�Js�Jz@�cn�R�x�q{<M���@���y��{�vݪu!�B]�����ZL#B`�m��`3�t���![��H��,��
����ļX7�r�E��z]=$��,M���&���������ʴ�"T�՗��-�#Ųh+��mjĺ�j��*�����m�U�"�g�\,�nҾ폹�+�m|dK�M?6��en�wv��I[�����^��>6%�����o ~���*��S=��U�����XB�Pb�q��,c�1�ғt��ߐcnf�c�^m��K���ąϣ��,0G��\�X%�Mn�*�Kq6�F���e�fd%GȴF��Cm��]�,���
�؎�4����U�t�xoT��\��:{�MT�L��ˋ)F��G�k�u��-�͐��2-����ɿ���h�kU���)�����'��	ٟ%9i��I�I�V����Kd�$�˫���ڒ)��;z�q��~��+v���W@f�!���vꘃ����K�-��AnJ03�+������. ���'���to�`EYΜg����Qz�G�� ��ɬ'�U݅�� ��O�ӛ�r��Ҍi��<�c���B��k�!�#t�ߋڤ�5jͣQ�1�Z4	���L�αxɴ45.����~/��E�|�F?H#��H��_�M�`�ۮ�>�H\6��U8\�N�(Yc ��@ʊ��;ߚc�,FZ��Y×�3�(;K�f�V�V�s\l�(�x�R�-�@��d�6�"�%�^X7��/��P�ؾ4�R6@�=�*����~�lsР��qL��d�ܒzs.S �bh�L�)I���?�/i�S�ٽhi5��(��ڟ�,�«P7zR�3ȇt��hg�fk>~�)�'|R��|{&%�YW�$q�5�r���q�Âc�L��A�J`������	�!����CE�7��<c��b��*�KRWE�ć�b����x��,�Д
[��u]Ůn�9��h�/w�"��0\�U6�`"�}&n��bc[�ץ\\C�h��J���~t�/�`D�fEF��YP�df���W>y��x�i�t��<ڏ\P%���
�i")9�i{��C��󺻥Ck����8�"`�j�2~N�e�Uh��NmQ@����k�E�#pQ�Kl��۱j��y�*�%cJ��GX7�^���}sg�X��?������d��-�y�}��5Kw���S2���rOHKʻ�Ys�"�}�G�����mx�����������mk�r�� �-1�c�鿆�D�A	w`$�R����0�沷@�y�e����\OMp��������W�w�L�m˖��R�( gI�43.ԙ>%�x��bpc�a\�G��=׮��ǝ�;,ns���aY��2���s�SU�z�|>�������E2��i=�X���9�k��FKA���ƾ�3���/vɵ-A�� �����D���d��J���{����޻#@)Dn��$Y���5#�3����@{�@�L���}4�H�	�A�(p[��G�'mu��5E����q�a�%&�:���m��֔����Ћ!�t�>Wƪ�E��k-h������Ͼq�
���P���`�+�L5g�L�WOo�ܰ���@��M�Q�E�NLyX#���Ao[�-&P�H�̎U��PP�_�н�c�����߭sp~R�y�4x��?%��%��� �G?��h�b��I���/q�Ԅ�z�	�o8� ���pt�����G"��t��%�ŇєMl9g
G���E���M��p(�͏���a�%��������4:�O���qq�r5J�T�ZH�u�K�-r��U.J:�|�M�_C@e*�!��$d,�/Z&_�☃�σ�� ��?ev�vz�Z1hR2�|_��63��Sm��\VU#��A砟��`����� �s���:������ �񜘳��"�X�#���`�Y��Ѱ�/�%J+/]���@�4��ނ�.w��$@0_�ptY���Q/��ZsU������	�;[I���q��r�c���oI���׮UTT5<m��@d��V�I _Qo�2�#Fy�mz{����<�M���~�u���ףunho 2ۨԯ�xS��'�I�'{�]�>^RJĽg�&�e~f������L�5h��|�PK{�vK���I�(<~��_$�!�e�0��`��v�*
}")Y�Z���h��џ�w�
���M��Z��jnyt���8}y��%�Q��O�Ź�g}b��1�2(��j�c�>�cȁ朜�q�'��?�����(�)R�F��Tt@�?���?⮟�NC�1�2����m��o8+����NVn��3Qb�DD3Dً�v,�u��@�@��w�-�h�k�l|�_J��߀5�0jk8i��A��lT�z�*�fM~��4�&�qM)7�ή#�w7'�`f5E�Z!��%�|�-ZI7��m!�@B����v�d�rP�/�7� yfW��Q~�ml�
3wR���f�������-{�h�p@�a����e�9]�nfTޡ�n5Q���l�)~�ϕ!�>S��$x�ņ;~~��a]m���t	�"D�q9Zv���?�����N'y� �p�r�g�e�|�MO�2�J�mq���ƫZ �w6BZ/xZ�߲��o@���й}L�U���w���j�ps�U�Y�`�X�M<;i�p}VЕv���?W@�E_>�~9��e��kѰ���5u\�o)Pd��LG��㝝�j��%2�Kf�"=��~��P���ڌ�0sdmS�D���`f����{�#VCpV�.�Bk����`��q�:�܂'��7+yz�F�"�+X��4W��u�����s'��s>6q.�+!�^��gx3�j�>�fϑ�ѧZ��Q���k!}!މ�����Oi�@�F�O3ZsOgK�R�5oR���W�X��U%_mi:�%2M.�H��Q��o�o\�U�X��H�@���j��F��@] p+�ŋH�rj0�-hn��K��GO�b��"�ޫ�y�D��4������6�`���:IH��B�E��J������Ś�A��S8�@�`��5%�f�9�E�厸,B����}T[�b�˭*���#���S��{���oO>�>��'ݩn�jG��@w����KL�iƣ\�ؐ��~{��>�����B�8��?�G�	5l�&�����N�*��g��L��J5&�=Ӆ?������I4T
��a<&w����� ��z3 ���*M+z�-2��=M7��_��!nh�{L�(Æǟ����=���YX	�LxlkV?�N�R����8�$������t*E nthd�k��(�vb~V��(w1��i���"I�q�:;g�h�
����"�����`��K��C���,�:���u�i� ��s?*�{�x�k.(���$zE�!�����~BT[��\Wpqɥ�B�c�1k�C��#%4�۔��"�C���u�v�?Ol&H�a��:{����_�l��ю����QI*\GV1+��y}W�b_T�ZϘ߯DR�\�Q�fQ86M��N��T-,�.�(yT3�f�=B��W�`5�(X�XP�2v��W&���*�_ ��.t��0�a�@�m]��Kn��V/h���U�'U?�I2�]_�@F�Fj٦����ҖIA���-�,�<�45K��q���t]�oM�����G��q�ս(*Lף���0���?ma"w�i����=3cH��}�[0Pa�1�%Z�U�:O	~�(c�����a���5?˛��S\2��i��~=la\;��Η���k�Ͽ+�*��O�W�'��#n� ۱9���! <Q�o	�v|p��,�9�j�����F������Q�C�,��[���E?-�R�q0�e����u��J�I��8��ų�{t�с��d�C,����� zq�NE��U�˶��Qy���0]�'��}�-�¤��L�l�i���7ұa���+9y^9�N�>q�?1t��xǵ�����C�U����͉�!���O��#.���^�w"q����+']���[[^�(ҹ?bcK�����R��1��J�������c����x��lRO'$+�&=��H�`����gw;|3IY��~���gce��hE{ܤA_q\���7R~DE(!�x�a�j��J�e�, u�s[}d�.$T��2F*:Ui��>�X���PD}O��YG��pR����tC�>�Bӌ0��-,Z�"�tȆ;d�M̎F���?��_T�$�Jg�o!c�"�D�A�Kb�*m�5An�����rӗ����E�-Jt;C�X�_ԃ]:��Pʬ����R����s`u�'eK����Y�X�m~��U�
�y�3�4(�����}�"�|Q��Ȧ���:Df`\"�	R)����b]�/�/-N�@��)����ܰ�ie�5<��d��֫w�n�q�Ey�/̝摹8?J/��|!������+o2��r/­İ~�-y ��TC��\Ѳhj��X��w���^ڜ�U̠�"��t����>u��G�ˈ\,z�h��ti?"C� �=�3�F��l�<��mW�hŐ�\%�!S�b<!$��ѷ4�H(��TM����Nw�˔X���]db����^��y�j��m���ƌ�(��- 4�'��m(�� ��g�ϩU���W4%��^�]C�f�~+�'��T8�e�^�!��2)KUB*�`���c&,�4��f+ݎ,�����h��3Jos�M~LeV���_]BKwkUL�K:��L�J���	�Ų�g[��m��X�ⱨw�u:&������3A]h��䵨3�:H�t��9�c�/����q^΁�NU���Ё$ﹰ8őM�r�v�S۳����ɲ��S���Rc(+�	 �H�w���+�~�iO|c�n	��5�d�7&]U�ę�K^ް,,����p�GZ奷�^�d������5������%��� ݕQ���*��O��*ġ~��<������<��>P�ӯK�$OQ��@naHw��F��C�VZ%�[���X���צ�`E