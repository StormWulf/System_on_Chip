XlxV64EB    3361     ce0�T(X<ӣ���J@�����Y*��������V�(���$jg�\���_O�Ҵ_����z�ϸV��aN��C��g�8T޵�R6���|��|�0}"F�-A>D�EѬ$UֹݚH�+sbw��c���.�
;1��{I\ܿ0׶Ok��(!��6b�,NO���f�ّ ��ƽ}h
id��"�u ���cSd�MVi53�h�X���,���@}G�_b��>|z�!����7�x4y`S��z�;��� x�#*-L���Tb#�S��+WT�oB:�Q'��dH�����s�B/J+��&�56�E��y@r�o��en������n��I����.��T�̅�	'�rʝ"ω#�[��� �h����޶H� �.�=�2te�=�41ԝ�'������˚��D���/t�e�G���j5�#uS�Q��Tzw��mN��(�AT��;ܴ�z�n��$Z$?p��/z%1C<�|.++���4	�����i�eh��<������Ќ�e�NBVΗ;)6�G�\EΚ��|���q�L��d���?)4޼e�Z�tS����4�&�	�h�X���a��}(9��#����>��>X�1Y��>Ae����j��3��{La�n!o�n|'�+���`B�v��ҋ�j=~K�q�[@Aay���%ಕ�"@��B+*?��YO,��'x�>�����ѤT[C� $vx�U-��^W�$�9<A���!5�6	r�������[�ͼ�#n<X]����۾�z�\����pCB��'[@�0��EJG��9[��ΎE2՝�ށx�J+�v�n�5vc6�c�@�{X`�h��<-zZ��mˉ��l��a�/����HC��v�9�������_���ʘ_ɴ��mT�d3*��g��/��ͼ@I�I�T}�����^�_���M0e:^7l3�r����n�ۙ���
�W�k;8GȢ��o�7��k�٫�.��}�����"�§GwQh��%hr����Y��V���HD�	��=�^�!�
���81T#��QƢxxb�VMU�T�n�&������c��4Q�7���-�y�zÔ7�-�����T ���|���㕪��T
��6��a?G�k���煷	��5+#V`f��h*�:�$��ܵ�&��@��x4?�
��?��s�J�r�|`l8�W%?�*6�%��gI��;���f&2>��A7�M��Bڣ���"�h�M��bH��]!d&kE߾3
�XKP�)�a��i��6ufM�P2O��M�i:0�A-���LP4=����<v�5��y�=ZSִ%`A#���	��]�Q���%q�N4�ˋ`�%H��1"��<�!JD2`���ͧ�z��L^�	#�2u���b�,��*�s���_�3���r�y�Ѿ�4
m�+Lf�wp%H؟��OP��+�֖���i�wy(�i��_
G����2]�Ną]����gW�oU뀝H3�G g.�LQ��r_Ŝf._E`YL�7��q�f�Nڀ��b�7Y܋���EnQ5$(��um������V�u��Vx>�K����au	ƙ
eˇ¿�w��U��'z`$�q؞ڬO=���4�����/a<oG���b�6]���)��	Z#��tDFX-�3�y�zEgi�ՙ��5����۳��L�X�R�����H�^1�g�Gw��N�N��hh�B�xGY���)5d��S����+�lw|��Vp�lv_��yu�Y�g��:1(	Y<H��j˺O��-qj(=lk�"R49�T��D$|��=n�YWxl@��U�9Y�E��&2\��c�䴲o����d�Z��v�Y�p ��(�X�EVL����=�M8����|(d�=vQ�=ǩ4��Ṁ�X�,���e����1O���z�{�aƞ�ޤ��Wo�p���t�'"�e�7\�j�m��v͎��S}5l��O7 '� R��f��*��3c���C�UL������1���I��{¥�Ӵ��՞sb���5(F�\���nP�B�3�+d���Ǵ1�O8�^X�|���!�7��q+����Q��-s����n�~g��q�C�Eh���ٞIZQ:��V�r�U�S�lø]�����؈�|���� @���X�8z�R�b��N~Go�`M�	ܭ�#�7<+~ta~>��v�<�:��ṐL�;'������ʂ���cɽ��s�+i�=�����W�!$�j��/sƆ�ԏH��9��yd�NǄ���ۚ���\���\��r!y��.S�� ͤ,7�V'�	I��|(h���ˈ�g�yw̹�����l�>'�+����To�wBxiQl�,0;
�o���Gk�����Gj��i�'_��� 9��#h.��lf��h8��[����A����"��Dt�� ���%�t^�} ��?���V��:H�d�Q ;����'��
�p��p���/V��8����]��a��$��]4��4��pj�l�2L4`�X��]8�`�{��e^'�0�I#���ދ �Ԃ��F���ڧ'Lo�_4��w�#x|X�х�K�噁��(A�u�P�V�=9��Ÿ>lW�6�: O*M�����b�ƺ*����M��S����W [��V50���2��]�5��ڃ��]�xxn�<�Dׅ�G�k�>"ir� F����#�y'^�dE���6o�2��s`�F�T[iK�\� ���"e���Ԉ�T&c@������&8������jd����S	8�Y7����P�(ҝ��7�u�Y[�$w�l��v�>���J�����]"r�&�{J���ǖ��I@O��7���:cű���q1������A��_�V���8����� Er���.c�T���.���*�1���ʎFL�ێVO��Yq�7��*lԓ��
�=;�3藟$���uaG�)a���T*I�#�.����a:/�.@5�=�ityY}�7�'M3�gѴ^D#s�g��<�� ���N3FhѲ���LU}��ͻH�N�-R�@T=�x}�#�DX+�2|k9�~;�퓒G]���q���f�'�+2��HIVf���Ⱥ}��dPE�E�k�Fһ"���_�:ŇX)B-).� H���8$�lC{����%E�9T�M@�P�M{��C�Fҽ�j�T��^O?1���tiQ�r)�wc�GUSF7�����{�Weى�q��G�f�� ��p)K�^	�%n!2^FZh��������C�Z���87��dC��()�_�Hv4��Ͱ��oiwbp�3G��9�䴸�R�