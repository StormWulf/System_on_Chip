XlxV64EB    1b6b     9c05��R�=H���@��_�5�	g�qݳw�Ǻ���-��;{Ux�3�@���_7��5!ۀ~�4�t௜tc	f�y4���q��
� �� ���1�����>�j�f�0D�{J�@����r>�"�B�[?VC��l�c����!=5b�}TF��˅1W.�w:��{Nؕ�k;�6��YJ�Ziy6�֧R"��S���ʲ���V���6䟞�+����H8T��(��h5@֚�ͥ%�f�2i��=E�_T�r�2�r�ɲ7+	�]�$�߶[��Ok�ONaU�__�q�'ښ!0{� ��ױ��M�������������e6~���;���	����yL�|&=�4�S1r�BӾ�q��:�B����!�;w˨�7O��j����*�9#<���*�E$v	i�Oc��z-!��'�r�|�ҢB�y�ú��WG#ע�w����&�}	�\�Y�ڼ�� >�d,��3d���l̃�xd"Z�����KH��K�=vm���4Y<Q���r`�(K�P�E}�@�V��k��7?Gc��%��qS*�&�T�gZx�L'5�2�����B)|q;I�{�:�)�N�jDyN�?"M��fneA2��ja���Dl� x��x)�7��]L�Cw^�63�J�O1�]D�&��z^�m��Ʊ�H�a�TدD�������#���j�n%�ڸ
 �# �B*�]�tڋ�'7��#.�т\X9����q� ?�Xn�!��a�����$��T�6�es:��������^└�J;`�t�&��l��f�ej�CÖ��j�y
� zs�O��q���Z��ag�Q,�l�<�8�
��Ek��d���[���lP���|��P�/9�/8�i��I�̈��Nv�
z�����t�2]���g)Rz�+�q�֓F7����e�3Ǘc���=�#�E��:�6GqD��|f�cxL�_ܖ��?�����ir�f1U�����H`�ζP����{���cg�Q��n�l�&���wI���} 4��$���HWq�+OmN�P68zs�F˖5���-`�dDۇv.�z�pܩ�"�ߜ�M i�W�����M�$�5a���ƭ�ԯ��<mX�~ʩ׃��>_6G?�K�>�
F����fl�m�X��5�T��3�c��9��N߃�E5%b@�cS�玆�
Ng
�J�����{:�pT�����}歘���?X�}t����/�n!5m�V��.�HL�&`���59��0�N�*��?Rހf��W���ꛊ~�����U� 	Q�C�B�l���n��1�_�gHU��Ӣ/9)�*�&�<F=�m���TU��c��$H�8��$��x�q"��T�m�1�g2A|UNS�ǯ���7rbhꤷ�|�gQxT٤p�B6{�['���<��Z��S!�����d�,!�2�QA˶��~-�D� ����?������I�N�\��+��B|�!��1bKpNs���;'F!���A�W����r�'�eP��'�T�?�[������}�E��eGaV�Sݘ�tD��b��V[�a���U�+��l[Gah��������U��#h��^�7L<�o+-�T��s�rf���1H�n�5>�I��Z����%xֿ;(�⠅��ު�A_U5��z���8%#\�i�G�L�x��	��9..���l+�����Pλ�'�{��x��'��޸s�+�W¯c�B|?�lC(_BmmBI�aP4�U°��6]G.�k��6qW�Ua���⾇e�����#z�iEqx����;^+ǚd��,�F���O]&�{����rM�:eɪ��o�x�Q����9:Wq�Oqe�,��F��i���4��3ޯ0uIۘ�D��D���?.��B[2E���Y��7H;_�g�i�P�$�FD]�p`O��dĽsm�.�!��>�.WCW���F�L퀍�������������y�4�X�z��ˀfx��� /.�:5�4���pd�f�cꆷnY�P�J�yH��Do���/��S,%��|���D�����u�y�GY�Fr��q"	�WQ��FG#����El%P6FD�h�knR������U8�ԋ�g��6i�Q?<g�yw��,��]�>ԣ���Zh�)�����(�gi6N��WЕ ,;�X_��im�]��J_�r�+YU���pO��>��(�������@ݘ��ifG��$�0O��Fl�J���V#28�V����>�B���-�ΦS�,yon>�����Gy~*̕
. 8*���Ϫ�IeGCR��&�T�Yn~@`��9U�`ڶ�@��B�xQd!�@�*)g�?�!p�I�M� ��z-��;�U2c�U�}���s���}�~0X�0�(�t���9�i9̕cNw��\Z�j�!���Qe�?կF]%�x:�Ϸc����ґ�@鯨A7N��~xd���<��F����Q����(1G