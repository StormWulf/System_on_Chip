XlxV64EB    fa00    2c20��q�����Zwf~fD���	�t���(�1����E��A��}�Œ���{6k�x�vj3=Zn��W1E�,dĭ43d������뮕����ð���4��#�XVU���^F<v��B.��\(WԄ���_C�N�"�b���_xA�4)>Q��ѕ�U|p�.���m�`���� 9U1s���k��:��V������ﾆi�ԻW%���`�vc�f�ŭ��ԅ:ŮXT��)h;�J �a/C��C���_}LOz47%ф�������Iv%��z6x*���r)a��T^�6Z�`v�%J�J詅M���S���l�wץ����t.�#)��6PD�loTՋ��?�bd��+MFӷ$�WF<���6'��3�S�K')�ђ�2����mkdGH[�g�Ám���H��(4�.��+3��2鿑�q��&��Uk�<R���V�F� ?x7�	�<���=��9���w������Ȏ,�G��=�%1$�=%>vE���������ߑ�B}:�wiD�+r�"ʭBP�� /�a,�;�]|�M�Z�?9^wIS�2��Sg�#wg���r��0�O����}���+��9�5�C M_���ҷCL�D���n#���6@���[�u�T���"�0;���~�Ӣ�K&WŤ�ֳ��W(����d1R��T.��6IG{�P��z|e��K�����C����.Z������\o���4���M@x%�7��A@�tc�O�����3l�`_��RYә$;�qj��:Cz�{��G�K鳒���b1��t�G�!��Y㑣Dzؠ��j��b��,�;f@��]������x�a�ף���2��XK�S~ڵr3z�L_Vv�9��-m&*�b3Q�|&�A9x�T��	�VL����m�k��В[D&q9W��nwhJ9يŭKT�/Ɯ�(�S�T_�ֈY������m��{ހ���w�0|�$�!z�I\Xm=�=Ua?Ɗ0��o��Lp`��b��� h0��
�M�_��'��|ut*e��	il���c���۞�}�O�.l��:d�!O��u弶�풽�)�������WcW�f�Q���B��.9���\�^�tXb��o,�{�aү�7Q�1D�|��3y
�������#�nsW0�D現1�,X��gU����3;m��T�ӥ���	C`]�Uot�ŮVz<�>��=�[�G�O%֎y&^�/,Cpg/��?�Dw�.e.#!i��:�An'�]�&��u����V��2bp�������U��[}�i��jb�HU@5uϳ	F����#-��|�/����x]2M ]럓�ō5Z�Z�mOU�8�s�lE�K�;۬%��+�5DV�~��d�������G�����U����)��?�N+��7��mqL"���12��#�qDŚAi&��ͱz��+�B���s�K���b����߻ќ�γ�������^� �_�j��RO]V�����"��W3��3��0=�ǉW9h�ɓ�Nv���Ԝ�i}�F���U�$c˰Pٚ>�
dtB��3=����Al{a,f�Be��T��%�T�V˰dN(�4(4A�Zc�D9d8#��BE��x�[ e��|�V�p\�SUd��
�Iɞ|���A7aB�Y���+������
���d��A���Bѡ���K�^]��[��E���zÝX��""��ЈZ���7&J<{�m��f�(�Q�����M ����%l�ؔ&���&<$۞�E!�a���2���L��N��Xl{5�+h��&	��ʿE4��{.�$�F�c-j�N�FIu����#�e+�4���kv��9G�<�C��l��w�4u�3�Z_'Y(YY)���dO�x�-[?���!>YX:$���&z��1�����:���-�0OY.6m��l���$���0�yq8��#(��^�� ��7{ö��]3"�e��H��	/M��3掩�]2�J���u� �@��@+4F�mP�_��l1[(���fM���$�SR�aC_b��YU�I���e�ߏ��� ���L��(�Ϋ�iF��뷪�ug�����|�FҮ0�v1�{��y8�4n�U�	���'�#�Cs�.>�A�-`��(V(;�`��^�02����韶gƩ�2*�r�|4�~��?/�3�T��hW\R`J*��59S��e�)7`W���>���R�y�C��O:8�(�J8(�_�@����5�L'y`m3��Q���[�*��$7�%�\5p/��,g���A�R_W<�{������
�:�R���x��
'|u�PE�?
o�V9�����ݦ������+�D���>�KD͐�L,��D�����_)r�)?�l�\�:����7w��2h�ݡE����U66���������X��и�A�u��Je��!��fr5v��k������j�R�4���UT�w����H�����_���<�@�P�:�̾�x�h�J�p�R ����Ý�:��{S�. �ȷ��P��P�Wy���pS�^�S����Fr���n۩����%�W��b�"cWҴ�����6���7j�������B=?؉�>bxV5�C�-��f�Q�b ž;��U������k��+�&y�`�z q��ޫ�#zX��O����X���T�0����)K�]�i`!�a�)\e}ЉN ��߭i��O�� M8+[��6*/v�tc$��Do��"k��)���M�P*D���^,�L���6L�
[�#���&�	�q@:�#v�.� �M��
>k�(&I�ق��0)�ͺ:|/�����H��yH[-��oU\H]m��se �<G���zu�+̨�K�S��t�r�Sg�f�O�2���y@,-�#�����}��W�H���:�����ȟb��	?*�u^��+RN�)�XC�-�3T��lW)�}R���S�Ӝ�X���k��������Q�,��;(ˍX��6�
����[@;A7J�[Ԟ��K���9Ĩ�_��E���W� ��D�aƼ���Ѡ��C����q�40U�k��TKV�f|bf�hEy:����&��iE���1~U)���{��R�2~R�NEs.#�I�ȳK�����y�\���%��10Ҷ�!l�'H�OԔ5ǡ��yld��GhI��y��ĨsFju_�ȅs���%�ۻ!��OA $���P0=[(�g9�q�S�����U��DȀnC��]m�;����V�c$�E��������N3kp��z]��Cp�o�HUt��E)'�#� ���nog���d<e7;d������=�
Άb�/>�\���mX�������G�}�z�؎��W�D>T���ǓcR!������3y�Y�)L�yk��L�� ,�k˲.�s�|j��D���]Գ�.�,��h�VC�n�C�M6%[G �����3:k����f\�>��0���ьw�<<�ݏ�7	
��N7�'�h�ٟ���So{�n���l�KC�`��N+�=�6�u�2����,bT�9]k�J�����D́�~��˓X5A\�I�u�3MLX&������_���_�1�w}�dBC迈�.�ߏ�c#Vˡd�p�؀1�0�%�}_�W�-@T`�))ۣn�k�jƣt`���ײ����nN[��Q�R#�v�ٻi�/��7�Y�*��(x�)n׆j3@~A���Xz�L��f�����L����8<猤s(���:6����|�"������D��Qm#�9�)������&>B��b�-P$����n���Q�@��k���=�3���Tٜ	8���>{뱘������'�8�Ƨ��~���v��a
��.)mr�}���Ǔ��Z�� �j� �4R7���"��>pyUO���b����~p��q��va���G��Ͻc����o� ԝC�E���4B|<��D��h����BНe��/��}\?]H<��4F�ǃN��V�ܗÃo�B}I~o(�a}IJ���<RMã\��S�)�ڻ�M�2TעS��1�����ƙ��?
��z�`�?ͦ����kO�?<�͌���~�ꢄ��e1���cg�����1�`��޷��Sd��C����ya�!V���C<����t��Sl��;�=���sB�|��ED�:㱣��wio�L�	]쳒��C*�죔hvсcgW�#;M�[@,z�4Ĵ7����Q�����+Î��N��V5J��41�� a*~h꓄݉�E+������԰��}D����o~�ݲv�d��۞�@4j�w�7P�J;SL*�"�}VhB��<)-8Ҵk���]u�c]/'r�珁䠀dp񾏇����h�=^��2ڥ�kZ#�$�-R�d�K��_�fs�|����_"Ko�ٛ�A����q�:�$��qo�F9ɩ�;���U]\n8��'w��7˞�*T�Ӝ�V�5��91�ڷ�4�P��aחo?3�{�����Y7B��슀9Ϗ�.Z����|]|8�A�4�M����/�;�Af��▤��M������`���)����������?��9h�b�]�+�-X����ZI��i�Fqf����l���ˬ�w%���\S�����9V�$�U�Nh~���z�bڸ!{96	p���߷�vw����@$�A�M����e�-�@ ���T���+H=��2�@���g�4�p�N�4u�qV�3~���tb5���ʪ�0����e��u<r�c�ֱ)z>�����s����T��G�6�����泀A�R����wϝ{�g��[����/~ϴ�6��b������o-;�����#��=��UQ�\;�I�'v}>���Gɬ{��n��5�M���^���g�A	��5��H�t���R�p��l�% ܩ�ǋ�����[��{'��;!��#N���1�p����0�q3��m���3!�\��%�?�F�҇�z���K)6�~�GnW�j�9�6{�+A�!�G�q)%¾\��<��f�P�����P���.�'b�C&;�xu��o�����Ce=Y��<��@����ː��L�]w�����c��ӻ�i�h���Y��r��^w|Nsj�{�KF�f�1�4l�[^��DC� ZI�3�f�	8-S�nH�𴣡���e�p�H���jsC���,H-��W
�?�IĄ����˗�V��E��}�(L���v�fB�6%Bȶ�Fb�,%jU�7�\��0_�Ȼ&G�)[��ec�>��:c��:�V��		2r��?�ѭn3��A��/��J�����{Y���FcU�{�"D@A�' q
{%rsԘ�����ԕ{Œ����:AGrgkV[�L8�5�=�1Tw�ݒ�_w���2��akP"9 . ���m�P����ʲ���W�x��y�w���I艘b�����yN���_���Y�e�S���B��eMw�Y
.���:�@�߲�j��̷-���lr�z�1H
���� a3���/���\��)�M)�k�k��Kn���Θ�)�&�iƃ3=9�+��]�~��
.R/�	{�:>}:RE慐�%������~T��G[�$�)Z�{8�*v/���}�""�k|� #�LZ�x�/��pn�?�H��,/"z����d���6.Y�j�B���-�E�%��}��M۳�f�ʹR�M���w�
n�tpY ��G{3阏�L'=O��yy$B�����Ҷk�*�N���N���f���/��:H��2'�����ő�^��������B�6��R�}o�W��vo:W
�R\�~?��N7^�kO?���Ė���������nU�-����aQ�eЌ���N�=k�� �tA��Dz5� �4�����6�q��k�̃~�X Jrlş���rar�f9^�>��&^�X��/L'��ڼ%y�`v��Jz�9���}w����s-��W��n"s���p3u��n�������9*����^=���Ο�6Pc�@�|%�r$|��۪k,,`�XK�J��PesԬ���R��V�]���t��1��p�Ƥ�����⦤tc��V~�3�ԺS�	�Ws��v��~^k �Sf����u~�������@6��"��rB��������5<,s�I?'��$��A~uJ��8%�c~�:�8�	�ݛ񗿯�����Xiƍ������ov����,���?��v		��"��	��0�b0��ʼ��.���Y�(���������&�:�Z �pگ�/?�0�|�S%ʆz�}m��ܥ��4W#�K�q�,?]q������&P��91�W��^��CG<�/� fx�P�۲�y�������i/����4d:ss�) �����)��a��!K�������o�eoS�&��gJvf"� ]"�.X�f.��8�2��PcUtQi"!MOѼ�w���ߥ��d�I�^�H5�)��t��H�Y���C
#��% �k;J�
�!���v핌�Wwη洇ΙS	�k�OCd�+�b����vÉP��5d��������ܗ^(��T����3�4S�-�Vä5B|E��>DjsVu��t�ː��O&i�1��.E�1X�`�ƎU)���cL�M�N��"#�*nNu�&�۵s@�k�B�ຳ���$�~O�%�O4�kf[$�7���)�+�+�w��1��S����@E�gg�<̡�<��\
��8��>�70F_��6��X0�9[���QC!�&(�m6#�@׵Z�/������0C���Q��w���R#N���7I���I!�^�:�p�=nQ�v	�p���O�X��B�+6;���{����ݬ�Ȇ��^��na��J������k���#�у��2'>҂�EΧ�:�'8���o��mM9������_p�s���oI���
�~�-�2<bK�����אnȦ�+ZY�����z:8�v���7)�C㺣�aϰr�*Q�\�t�ܰd��/��Z�3���Weˈ6Y*!(�>�bz�(����v��g�~�F0�+)��W���ʃ��>2k����؁$�rB'my��g�ܓyn�"I�2g|�Gc�͠�-���6K�gmHz^vt"�+(1�M	5�elu0�t�C�s�lw����2���{�H7!
������<����k�iV"�S| �C99~���]K��cі�o*I���b��ᣟ�%sb�1i�瘥'D�^^��ZZ:����I"��(�����Ɯ��R��"�@<���-=%p��ԋK�c �H�wT�̞��pb��^�rI3+�R�(�;J�I�����d$�=$��l�P+������6
O����� ���uIό�iC�B��q|�g~$A�F�����udڼ����"���]���QB�������`Ivh��^9�ܙ��d*j���sޙɃ��PATZ�P�
��ݣ8|K��F�)/N��~7��8�+d�|놖���d�]��b藳U�"(\C;ab�着\�|K7N����Y�C�)���@����3��Y�T6ʤ����p�<�2�kN/�Ao'����2���X`�41�fuF7�� �	��)(-�*����n˞���?˃gє�d99��.	J�lYOs�ҥ�A���Z�e�����<^JM��|1Sn2wT�O�����)}zT�
c�1x�O��ho���i���R�p]�,#)/J�~�6;Y݆�"��pJE?���D��TXwO������z�W�<����H�m�#�,�*�� ������NadjņD�P���E\���6x��Ru���߶=��h,�t���a��%�+�q��@�\��>Mjфq�A"�h	h��%�����b���*Nl2Z�M~�f�;T9���9��H;~w'9I'�? 	<�)G��<̓�y�ezS���l�s�$����м1�%:t ��7{>mYڲ������ ���G����\ٸ��ܧ�]�����:�U�������a�)�o�
�j뉀6+%�+*65�H�'<���
 v�0��� ���n�{��d��"]48�|(W�]8@�)@�������v	#6T�"v��4��x3����Kۑ��|+V%ci:��!����НU♷-C��v�c�].W�<�G#1UL��FW�k�-	j[>�P��7yQ���S�t�	.�k�̥� ��"��_^��zv%�n5�jXd�lKx����E���M
2�6���`4bs=�w�"]�.��=��ӿ���܀�C��WO�ꂛP����CQ����ͺ��"�#^�y��AEp���9>�F�X5��@D?{�BNɯ<�5J��.�W��\�~JD��~�w7?�����(ޗ���0�G��� �#MYu�{��tH����"jܮ"%�|��@��-@��-s�~�vz��F[
����ȍ��,=s��$��,]Ԭ.U�D��BD�n�)�,~M��W�T���	��4�����}����43&��%,@���Y�b#֐&���x�������TaM>�,a���XT��9F�z��o��7:쌾�M�X�u�R���tt�C-nxm�&����TI��W�Q)ӺU9�1j�	' ����'<vR�	���z<��ژ����h��
�F0��Cr�"�	3�Xѓ� ����f���$����֜8NU��v�/zdH�a#8�=8x��O�)`�{M�
4�Q�x�]���j)a*[qn!-��l0�nc�gU�h�R�d@��'G��ɋP�'Gz��4��G�w8�R�\�94���i�"��e��n�!�tw�3���WȦ�D�������+�j�F���s5P�C�|`e҂�1&�,g�d2U�JZ].Z��~�$~��blt#�i�'��wٻy+� �ч�X1�[�Cgɂpԍ��g�Q��R���xfJuц��&�n����*��[Z#%����!��� �� ��#�w
b؍H�!�^���n��3�������~���"y�(�&55��80Hky�7�G����YK�˂�q����׮��Y��X�+�ꗑs	@+�����l�E��)�f������nt8�܇�s'�9�,;��g��K�M��V�_� ��>�&���*��ZeM�?���4L� [`� ���1���Tu��-��02(i�ΰ�W��C��w��D��%M�K���c�j��q{�����F��|�h��2�I����~������3�#[/��a�_�G-�8ʪ�5�j+�NX��S�����m��cK�# ��^�mȠ6r�J�N�b�ʳ�,	pţ�Pe�������/���,��:� ttO5ۚ�����X����FYô��.�i���bd�uV�;6&�׆�>Ȁ��3�H�Jf���U�8DׂS�7{#�(���y��G��'F�R�]�Ev߯��5�A�D0g��!�Lll ���M>g�?�ѵոu�������o�0�pu�-'�����Y?U�k�D�eܜw�G��s�����,�#[
� ��G!fr��ǧNo�r�|��_�n�){ej���X���K��j[F�t&����Vn��Q�|�$�O�A9&sQ��t{���'�� �7��D8*_"��N��ƚ�E���_-gĎ���]�t�{��ܴ"]�>�<��A|��y���OY�N韾S�qL�3N,��&=t�-!�4j7l�����a��h��I�|��a_��&	���y�9p�!bά58.Iǝ�(xBk�S�[��G���MJ��kK>�|��`��N��U:���4 ���(�T�78(Ȭ:����H��֤����@=Q���5�A�1ޝ��O1�O������d�r��8!6���� �<�筽$V �H�e-���R$��Q�ɤ�g����%՗zoQß���Jx�4ꪐe�W���� x�nIi�u�2ԸVlJp�u��o�l�W��B7��O�dv%���6����3{�7z��E�(�8kj7L�#��c��O��G�z ����ڕ �1����[#��b/�*�NM���+=Am"-D���]�\.9��C1���v��0��τ���g����o���� e�=��{f/� �j��qR��LcN��s\�s��%#�Μ���D����$*�Cq��K.<��ab���f,;Dq��{��]���Y��]����G�6[�S.��5�
�E7��B��I�p󶂓�zt��?�L��ehp���cZ��սߨ��\�i�E?�+��׼*�pV�^���7Q��_�k�`_�u{��Xh%f��E������I{�7��_�������h/?�x4W��t���q���tw��\�8b�{��+��أ�η�n�y�m�0�ւ���đ�ˀ�{��WboP�O[�(^�Y��bN�:��Ev�k��T��㤗���K�+�����a��!q��9��b 㬤Ǫ�����z<�}\�X�Mk�(
jz-,B�t	˘h��'i����;�����n���3��=;� +����P��'��{&%<�i��q���U�2s���t�s�N��z�l���!��֯��4y�#�&V|�+�����X��'�o��Xʘ�'S�yl��M
�����ٙ���Mg$ɶ4�m�NԺ?���hx�e�F֕�����x���{q)��r|e
�k�e�
G�Hq�n��f)k�Ή�HP�g���j�g,��:��cW��[����N����L_v}�0@���o���G	�2l���������!�Ѳr1����F;��bL|�L�d�/~�ZyB[���p6��,���U�0t�)t� m����_�F.9���OT6�1v��㩔��1����V������0�z�����6D
w�$�����)Y���ĬI�F�6W�­k��Qq��p2�o�&�����'��~��a�,'<H��+2�UـCI!��x��q.�bV�`�����ђzlm*z�����ň6&�FT�; �I�K���D8u��H.k�
�!��kWmQvz�r�q���sY������
QJp;�����H�Ҝ�X�QO�A6Ա�x��whC7~%������ܧ6 � �Vղ��΋ 	XlxV64EB     f8a     420�Y����  a�$̣H�o�Ћ����3��|+�æ(�nn^��+3��-#*��(LZB[���!���<P.��t���_�Y#�D�J@��)~do�P5�s�Kl���r[�D�'�Bf�T1�Ye��j2~��G����Eq�@%o���}�L������	�ټ��Ӕ]5��Y����#�������+�K������ic$T%�J�B��.����k����d���s}�����ܿ�����<��J��o����ׅ�vtݎ~�L�C0L�as3`�`��%��hW�T:��u#������� ��U�ϺFSx�'����լί�0���
y���|�m�X�7��zꃬ��+�[rr"n�nS�`l�&'<���Й�nԀ�Yk$��K����q��j
TŠ���s��	G�1��*�Xl�q�����yz^����ӗ<��)�Vg�;0N��dm��_h��U�T���Z�o_�8�H�+�)\���0s�,�&
R�~ƽ��qG���6�9H�t��$�^��M�yC��zGS����l�~�?�74B���Qu�ɇ�h��@k-��T�<+��xt���f�C/��J=�V�����g\Z�b*�:�5b�H��łH7��`�ܪ���(��_N{b3���s��⣰f�y�|�4��2ڕ	�_�P?)�md�2{2��RQ�y���]�<��N$�]v4�+�%�hɞp��)�-�ꃓP���)eVkw=��M4��K�<�����*�����Z��|��.���U+s�j��)G�Ғ�w�/}����$���%��R4ࠓ��sh�`
���g`Lz��~&o44,���/�
��>�,B��>12��҆K�Y3�$`A#g�;�~uØ����LS4��%7@�^�
{,g��S�8N5���4��M�WZXN�7a~u��	qr|���j�8匜�C��!��5�G?e�n5xi�����zC�\�T�OT\�~r�ƌx�!h:�b]���V��v�C�4Aʎ��5���=ֶ�V�_H�'E%��"N-W�����