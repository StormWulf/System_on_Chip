XlxV64EB    2d33     a80	�
Q��!��� Gʈ���7�Vk γA�B�u	��jO��A�3,i����5=���d ���;�ȿT�'�Ĉ�`�d�'���K/�A(�E�ox8U�~=�A��,r��օ?1��a�tW�2s�U�՚�j.f.�p.p�CE����Cm?�o�1V�P��3
��7f4�9X�i9r���d��A�� ֽMZ`���8��%�����usv%�T-~���*܍}��\�_9�WB�n�$NG��.]aB\ֻ��C�]��5�M#�5�b~3���)�-N����=��3�i��e�|K^:�Wf�CƼd�%��$f~iyTW�hZH�yl6Ԑ��D*yʭ���x¯˃o�ƣn����ʓ��T���y�У���2��0�Z��Z�Y��
�M�IYl���x:�՗2&&j��b
C*x;vW͟���:�#��ɍ���6r�H�V5x�C�|��3O��{��0a��GU �RRDB���i�:�|3�7��x Sȓ��o20\z<��f�r�E0#8]b�&ڼ���d��b��>���ŗN:�8�?,�Xy�?�K.�D8O��ޡ� QW�9t�����pΪ�N������	�lX
{��cS���F���� ̫ ������.�R�Bjx����"�Z�����Y.o1����a�s���p�%$�A=��,3�V�H׆32���XO��{�"�������Vv�I`[s�[�M7ϧ��t�a�9x-~c������_k��qJ�";�lBw�Tfq�����T*+��\-���(O���\��fNx�)�F��җN��!��ՔY��u��@�Bi-ek9&:�{�z%|l�ޱ�;�*'N1۴�1��aO�Ѕ��%`����H����uW�z��F�9�x���M!�e�
	j�1؝�h��2V���A����u�5K+,�,�fJ�av5�{���^ʦ��M{D�4C6~{:1����,�}���"2��FR#�1�!��G41����;�򼨊��s���2?��gSDG��zb��		��:d�Ӏ������ɑ}��Zq��+�zi�|c�e�":�Cղ����"�3�Ys�Ss�y��H�6�Juq������b婺�[�y�G�LU'N�^G`�͜�Y@�D7�6DH�P/|Is3��e���'	�`���"���ڒR��_ڃ8�c9nS!����3j	��ZmB�[3�!��8����r���OG��qJ�\6�wJ�����R�%L�Ii(�=~��RN�P�a��
O���]-?�(�׶����X���������[o���x��8�&��Iۡ`������~�~�7;S���I&�j��i��B+dO��I�ÉMQ����t�,�mj�kO�<7���,%��UD�`)�*�/9:�*�.��%����|lY�;��^?<z�g����Wb0)�� ��HPV�ޚ=�I�����l<�g�<��WT�P��c��g+�#,1���4���W��x�E�9�Aν��m��x�\�3�.q?S2�C&t>��4�Ñ�p}����E�^���ւ��i�b���#�l��^�� �����rn���>d1��Q�F%�_��.�Mp����Np�<�f_���$�5ҷo���`��^��v|ҳ�O���B���<���YV�N;_U�M6�1HUAJA��_�J��G��Ö`�ʖn�/;�m��J4�)��}��'��Ҭ�Z�VLPIgv(�'%��cJ��r|v�g��<��+ ���X�����:�|W�O��	��Xd*�Wct�r���j��Xӧ����u�ەz1f���]����*G��-�m�����/˦p��{/L��O*���RfHDQТÚ*��w3H7~�����E�{0�ɯ��#�')Ȅ�� ��,������
�Oqk'���������1�CZ4���[����{��?�ٽ���95�@ *x��#8���0%s-�|�e]��|��֖ل%���I\�Z]�����l��)P���E�ۃLQL?���ݿ��w���	�љ���&sLHQD�º��b��ܮ��|Ŋ���p\���Iwo�-�6:s�.DSo�/a�������[�����	b�����1~�f�&ObS�����@�X��$�Yʾr��4��8y�s��q�
�NXN��ލx�X_������Z^oz-���f"i�R��� ��i�h������U��v`�e}- ���$�}<�uRw��g?\�V�{��6���)�F@�<��J�V��������y���+�X����B�c�4T��m���_	�h��޼?"�n�u�0�S����0k8 �'� �/&��R-~C��l���R���ߥg��9���8\��c9��M�Pj�)*�I��n���pl�*8$�?�F;�+��}�R�&�}�u |A1���t�Q�f�_⋠�O�?���9��]�0=Q�m�����D���ֳ�>�����Ws��s�5�J�R��W$�n�"<g�n_�� �f�[�� ��s�D�&�	ZGN�T���g'[
1�C�{�^ݶ!�y+!ѷ4��l�0���MAF2�o7-0kȀ�o�&w����6�C�mӔ���R_����\�