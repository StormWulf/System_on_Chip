XlxV64EB    8a6f    1520V2z�|V�.+���#��Y�G@���hR[�E���<>o��H� �u� U�� '��c�ڬ��,���OK����k��S��;��}]�JUS|����43���[J=�0�J�

�,���W��5�b
D8��hʇ��۟P�v7�S��H����8�k.(���бD���=dS�A�mՀ���}��B�W�1G'[WL�\���*,������ޠQ�ղ�0y����2��*��$m�\���O�v"�����T��B���w��ߣ���"0�cjh�΅r�*D�!��?��w׵g�����6�o���x�L����aW��k}U={�l�
p���hA't�鿆$W�FJ��4|������~\7k+;��(
�c��6��$	�kO_��j�����>7ѧxsQ��Ӏ����0��%���ED5���
T�q�@�T��W�|��3ᶂ���o���v�섮��>M�� ��G���2~5�ߍ3F��f�ZkAZ�d`6(!�ŭp1��[��O 
ES�=���4��T�*{[�,5>f2���:!�}��Eb%�}�6�f�,�7���\m�E�_j�qf}��H�O�u
�I�3���!=�-�>V�u�a�����"(^\��XΏҴ�
�I�<�ӫ�9dn������"�:���F��0S��&h�~6�G
�#�iW�*w|���N#m�-��&��/�L^�J���>����ረ]g�1]7��:��hzH�=m�"[b@�U�����Ԛ�*�yE��w�=��w�-P|M%�I#�eY��A��_: ί[����ȥZ6jpq]�b�{_FѨ��ee�9����l�}7�N�����x��𘽏�S��v�m��
aOq#��E��әg>���XB��e$��S����:�YC����$�8��� 3"/`�?��*rG��j����Ę�v��� �2l��~B�g](R�Q"��nL`y�=. @²��
3Ҩ��F-�/����[a�y8V�-����1�r1p�G�J#^[:G��|�pZ��-F*���,H����R�	r$'��gR�I�j+�knȏh���rkZ��?�faJ��^|=kIl���th�jm/��nYIn�3X��숩�����^�7���	خc�>�O#����Q��~^g����
�=���ש싋H�P�������J��=N+)D�J�цE�!J&eFp�i9�z��Cޜv\�O8��2�Qw�׆0�g�ħ-�N>����>3�[������!�b���7*?�c�S;��?#�<}�ә7Y�iLX%/���Y͆wR���~E�x,�����|5_o�F�P�Wc��qN@ڋ������ӎ��'[�!��%�6�
����sjA#m.����=�C�Ċb}�\��
|a3t,E�׽>�:N����a���b[�0�����>�cl���ߡ�������ן�����L�:U�����$.Ytc�ƪeA������QdE|�(��� i_��S4 A��ߺj�{KoO9j /g��B�Y�Ju�&��x�P�FQ�	���Lv9T�*0���4�����x^�J��~�B��k�w��"��m�UZMV!�S��@|#l��P� h��G=`кyi#r�r|l&Ulv1�C��u�x�|r��^�E��A��x�U�/?�8�N��e�bP:�� Qo�>�-��¡���Q�V���S֘mQ��@����I�SWi`���G��X}��d�d�/}����6�6���Ȭ����_���t<^���
g�6��֜�X����s4Q���g�B��\�p�� ��rӁM�	��p�5ZKʁ�Q��i/����z�7��4q�&\ʰ�K��MQ�dUw�@QQ)���v~\O��!�0:'�u<I�K�G���آOǲ�vNK ���Pm�z�~����ww^!C�X�t@�j������`#M4l��?�܋F�����>��S���)o#����w'���G�H^O�t`(XB�aL����?�(��D��:#`P�i!�ׂ��P5����?�R�b���
Z-���` 2�i���"1S���C�����_�h��Ι8�O�ʶ�h5m@F;�^i���'x���!s�\��Y�z+���d��6�F�Ji�3U6ClD���B�(?g)o,Qi���)t��`��%*)]�¶5X���*Ag�����xs�D��0n�4]5��0�`��A�;�#�Q��1�)oH���J�e.�o�ӗ��ԣ�z��$��Q9�@�r����:o�F�%`f�)��C5�B"#3��U��
��̦��C�88Dl;SV����0�ҔoBh�<������5�D �ס���\��ݷ[���z֯R�L~���]U�]>2������$���j�W<����{���U}��rO�f���3uSŏ�@SQ=s�=J��D�3>�}��W���r����@��毮]EA �L^ɞ���ȟ'�ihNT�b]�ɨ�]� N�Z+���g:1z�t0����rqU�Ε���䄠LZ��������ӆ"zZ�7�����z�w<y~���q����Eb� W1z3�����jf�)�ƫ���������ln5�Q�UN���^�	�_?ՊX��k)a���E5t�����=ܽ"n��Y�ﲿ�ʯƚEt���'4By��$: v�7�o�BXg+pK��c�5�#��TN}m�ܧ�)�H����V�p�*�+b�֭ [�a�[��g/��!'� �	;;@+��g�#��S>��v�1�o�	l��w#��R�����G�<�9��ރ�?(��-��xWF><�z'���S�w�nuغOkaP���,F!zd���9<�X|5���K�^9�	�I7彩�k�+Q�މ�β�ez��7��ÌlH�gL�U�eE�(GR8���Kizg0㳱ˣ�(\Y,�#k���:Қ��^�F o��ؠxLꞇ*$P�����A�J�=����sIV��x�T<��+��@��O=>��?�˒��0:�����¾�"=	����~�&[o�����i������ xBv�Ff�6��.�f���Y��Q��{�r[��w5�4�3�`�VJ�D	BS������5}�F��n�
'� ɠ&{�������]�V6����Ds;�Wi���ڕ��^3%1#D�+�}2���
3���� 0ĺyz����/s��Cp)n��vk	WN8`����Ik>�0�>w���ΑN|cj���7
7�y��U�!�h�W�X��g�y����Yj[�CY����5ga��x�^�q�(��0|� 0�t�*
�V�E���\p�*�A��haʅPp�E�5B���p��:gR�bc�!�g��-�&<��5y�]yt����w	����l�֫0�� ����n6����3F�Os;���GX#��^��n�Sg�T���N�G��bZ-2AF�[2��6��w�4g�t��fo[f��-6>����~�Od�kaG��>.g�);η�=��zxGs��k���JZ�rp�+��bOk1V
L�T����=4^;���瘙���嬺����f� J��hS»�M���|SM�Y*��'�$Т��C[������0���3L ��\� �����fY&�ěIq��r�p%A#� ٞ����N.
1d�;ܙ75Ui���IrŒ�
h=���]���"{��A35�C�*P�9�-IE�X`�y�mx�>D9���}k��x6�-y��>�;&����x���F���;�q����R�L�c�{{WH�W ��G���Ƭ�\��m뵀o�u9m�os[�<Lg����_�rb���Dh�UPS5i�"�/�{g���u�k��^��\�g&\�%E	���������/%�-!\�v�/����h .���䗕���ײ�5
��Ø��B�	��K�$��^����	�� ��P���5���ع�M��}Ch�C;1�� �j��������ʶoar۰�˿��3�A�Y`�tB1��ɊL��SA{܈���=j��"�RQS�L4kut�O�b�}�*��ۙ�[�Ū/� %�]1�f�'pG��e�_��[o>bA�ײ�N�B9�w�gМ�]�K��0��e�Ӂ+G�	'j�;��V��`��n�&�Gڈ��+���lG��{ᩘ�oJ�G	�0k ��=��v�U_�ԻU((����DØ�-�Z�r'�٦m�XMB�~h�te}؋���&	A՜m*�Y�X��ǟѮ����CT�(=ޗSh�_���Z[�&NJʉr�
���'�:���T��X���d泌m����3z�[ap:	V{pX?�<�p]�,J��ڿ#�B>������O����� ����!�u|y��m�ۚ��Ɲ�@�'a�9���]v^�]�Ea�7+���x�It����5,���i5/Nu$V����|�K��4a P�R`��m��Na����Y�����u	/W�xiȢ2��e;3"B�e�����L��5~��KԶ��P=�Ϣ�Kr�@K�Ey�<U����g°�FQ ��m�)pua�='TGt��n�H��76�?Z��n��W�-���˯�/Ɲ�!~��uq�'Y;�,�ILqhFAI��E��y[��;��h`zXR�� �����R��v�B�l��:��)����,ʔdzJ}e�k�p�m/ʄ7��P0��}�'n��|ֿC��o�<f�xQ��ޅ���2�aJB?�����%(.ЂV�c�ms�y7Lj@�eJ�d��<	;k�p`Sl%����+��L�gچ��i�R�:#��q��Gĭ���!i��M��e�޴	�bvр>;M��\��<��'�s�ߙ�Ý���*nJ�	�o�7�90�_=_��
��]y�@��V_j(WdH�ͥ�J��s��y�*�)0Xյg�,$�"	fvq�[]nE�g9z���4(ZFƇU�r9��=���4np�, ��m���G�ԋ���?L��������g�K��2�O��=,�;��\�Yi���<v��,2����2��X ��:Z˱���������o���@��~<�'V��]�c��x�79G+EQ�/�k���,%J�J�6����8����ܳ�9|�8����rg�&Bs��i�ҿ;|�n���p�?�ߘ,�5N�uʝ�6�y$n�4���5�pkSpN�0lL	'�uSmEE�2��9�o����3` ?A��Wc�@<G��&��ҥ�&3�7� ��Ɋ��f�Uw�`DS��p�QZGC�8�(i�8��*@y2㧮�,�\	k��4spDyZE8oԋ�:��L3�`:�c�)ϯ�u�{2%�S���\����y�=�
�E�=d��ʟv�ݗ7��<�6���