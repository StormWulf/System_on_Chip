XlxV64EB    2c29     cc0YZpq?��ڑg�lD�׊>Ep��	�=��+ců�B���B�Y�kV�����qzG������R���>�;V����V-q"a�zv.ahx�I�Z�^�����]	�5�R};gl�JX�?ʣ�J6��G��݇�Z�
��,��-)l7�%�-��\��2)�:��]��4�����"E���L'�,+m��%� ���# B�\�-���(��A��v�Ed䨑8ڵ��O0T�I'�ɦFr�S��D�y4�!E����td�����Q?�o严���#���(�����OE��6�T�$nw"t��t��K	�NP��\���y��ǋz��Yz��L�y�T�	���gk���'*e}c��RǗ���	�`('�NU]�`���E�YX4/zA����X��p-��gDa�-i$j���^C��_����x����++
���I�\��_.c��t�L�+��8Ē~hR��4��1��2\e�N��i�A�o����߇QKق��A۵NۖȋA�e	��K~��.����a�ꁊ����|?��'s믮<����^e���\|�G���n��+��˯U�-�K�$�i={nH��� �wR���I�5��� ��Q�Y+.��$�-�eCώ s�;��o-;7�?2'Z#�����z�!di��ٛ]3^�&�b�9�_"C!��2a���@�p�����.�a]���Ní����_J�@��Y[ ���v�"k6�:J�� �);�s7/X<�����d2f��_��Z&�ڒz��[�s��q����_���q&��Jl�r$QN���Ϲ©H�f����}pF����<6���=]'�h�r�l����tj�]HA�v�rXJ�j4�Q�gm!�:&�`�Է��@����Ed��L��z���(d9���������aw�o��#E����/��N9#��mv�B1�#V�B=�߷�z\�±��[ɛ�_s$�I�l����u��C>�����82,�5�5T@ȫ�P���{@�� �w]�CCO,ՔG:�Z�̵�!i�=�>؂ڛ�
c	{/�?�ʿ��]ЁT������Z��2��%^[�ߞkzyv3<7�HM�V�y�'�	�4��׉��y�ł�R+��D��:�l�-w��� S P]�9b�J���.rB<XU�	�2�q�a���6|��Ȗ�(���^��ܿ�H1����:��zw�<����k̺�.�J)Uh^����)�a��N�b)ϫ���]35��%�s�ۆpҙ��hMqr��1:����e~q���R45`w%��0}C�h���e�yul 5]�O �z8�6�S����7������Q>��'�
?��	Z�4&�<H��*�/h�s��d#�e��4(p�_"J�#�g'�囓Z
��V���g�y&+�"Q�Sw�L\�(�p����C`��Pr�4�~ �B&�#4F�R���8�&�Kc�g�U��8|9�c�a;��dh-�����?Ev� Ъ��g\�ϛ�����q�Hj�q/B�?��;nܛ���.%��QoX�h}^D��1�Vg���U+�&���Ut>�՘~���A,a��~V�����t<����{S#��[m�[;[�.�⧹E���T/����1�å������A��|�}�G�I�@cH�>�B���� S��%^���b�mM{[��A[Vq���#X��9o��Y�Y��cٕ� B��/�vp+�"Gv J�&a��1{:8i]�L_��Abە����Za~ԪY��ޯUd�a�b�	�X�52�֜7.�R�*�wo���Tf��R�:1V�\W�uE{7Q�#�m3}���D��ɴa�F���NS�k��yu�b�y(U��=t�eH�cLH�NL�*d�:R��4�N�+���,�����pkOV�`�xX����\�� 8:��z:���j><90D�����;�@Io>&S�S�:�L�tf���Qedq���Ҭ`�U���+ 	q�-W��x�p��zP8�R.gr��0������,���|�~J��{��X�H�/ ��a���Ӫ?2��Bt�7U����o�Mo@�7���q�֏ah�b�9*�Hŧ���ߡ���Ay.׽Y�������U.�
�H�L�LC�[dy�b�����$f'��_�ܲ#~J���]����?/��3��j������TP)�>�3�ޤ�(�X�jF;8p�1�0w2���aG��O��2��d�=ٗ�z"��8j�z & ā]qp�q!j��-cA�/+���Ҥ୫��u��r��%��9��;��q�R��T����|�S����A�
��;�I�m�t#/��9�x�AM��Օ8����F�Ξ/(W	<1W6%lu�GH�]�)L�יnT)�ƻ��
dI�&U�nKa�,���r� ��mLE�`/{E�M���#�){JoIs=ڃ����~���[c����xk�j�ล����"
�bL���?�wiۦ1͔X�(���w`�8i��R�c	 �I��*�$��mvU97�
��z���/�l4b���<b��^5����n� ��XU���h+_I�쳐)봊ǕX>ǂ�ͧ��9�*]y�BӉ?т�>_t����,b�s�4GV�e���𗎥�&t�3r䄥Ø��nQUX^g�V�0�9YfDVB�u|�pj*/���n׈�����XT����(���a��)r��bg7
�e�D~:"p�#*�����諥s���M{��sN4�j,�(��Vԝ�����ٍ�e�ȏ��Ս��g�r��Y��H#n!�Vs��4u�;.L?��|$���w/��$[��>�²b�Y`G��t<��\Yc�dn�;���Cx�#��B�,� ������$��*���3��7�oG�[
0NA�˻�
	]7֝oT�R>xv��i�z�0�i}�v/g�6��>J�̀X��NX��>�rd� ���=*��4m���blM�K�7&Ʌ̱�_b�68)��u/I������NyL�7;W@D�6H��;��ފ�x�5�T���[.����+٧M��p�]��d�N�s�u�����&菄�p���~���~�n���-L�k'	�R�$_�v�7y|6sK�#YF1;�����bo*2�����~9~ې����OOl��et�U�y^����җ����Pz
j}���j}�����TxO`�lB0!� ��i�Q}�(O���̾5e �jQ��0�,���@���x��r�f�.