XlxV64EB    56c2    1340eT� q�#�X,b���/u /�����%��#�;b��2(��b�?]\�#������@�D֠��L:#�G�ICЇRs�Qw����b�^`swn8�}a��qq~��r��<2�ѝ$Aƅ����Iň����E��3B�o��*]�z���S���H�uT�7�d�0m����;n�y%>?�d�8>U��5w�B�[�ژ��C��4{���`z���y��_fV要�l�x�Ui���7XZr'Z=	�/j��� ��C�gp�4�=-y�<�S1[���_�A�����8(�.q6����1F�I�[�OE�jqtb��N�CSZOj��c#q�2~�J�g�����rg�?��Ռ�x�{�a=*��������$������`����ٿ�Z.pz�w���e%�2���q�D��8K����m������-QA�͛7��4�u�Mb�w��Rg�ͦ��'�:�uY`�{l��̩e�?�}��u:�|�:/��,j��q�*��-���C9�*��#��9� q/�PP}t���3��FS����|�Tmˉ����*S����( �<�CE������bʧ	|?�S �!��\w��\5Y)�"$���H�H�EOX}�����V��5��G�_���l�����*ܖ��m?�eU� �mu�'�E�>��K"X����_[�p�c�c
�^���CΛ)�G�������`��,t��fR��[��������1*l��8m���d�iW�3����v��b������ꪡ;�3��앩s�@�q����)�>J�>e�Ս��P������A��]8�4��)�*��t���l�͑�%G�Ƿ��]������2[ލ4���y�����B�������h!�Uwq��F�zX��y��G��/rQ��7Xo�9IЎ�<����W��0�G���/����Ѻ(xH��qJf�W���N�J�O4Q�V��!5��u�)T��t�Kޅ�O�֪���h��������m��`o	o/�n�JǞ��+���R��a���I!o)i���ei?�!Z]���<a�H~2t��f�&�'��8)g*��u*��h�o�G6��Ɵ;�S����f�-��6�br�)�o�ָ]o����$°d��:�{w�����(�D�ϒ����°���������T�����m��8�D_��kI:ZQ�i�9�
7� �8�e��(Q���Mp��q�V��=��}�;�F��i;ܘh���Vb*j
�o�]��P���HYl6E&XF��O^j����ny�Y��մ�Ę��jw���ܬ*�%�.]����hB�Q�� t"~�� ��؅��f��LOL��D�:� `�}v�O����j���;ܿh��.��F	��gu� ^rs�
KP`�lR4��P{�K�����<m�P��! h�؅�"����'���%��TZ^[P�*5_'��Ѕ�.&w/�QCAؑ#������g~��Ӗ��0�����s.>�=���}��u����)s�L�+��>R(�2������G�|���)*�%�'���>�E,�x7�a(q��D�����X���xZ�art�zU�ls�W��n�a���ථ���M5�]�J��׭��_���մшd��<�����Q�쪆�`.��bFhi��/�0��/Dw�ºF1���EPW�� �1u�t�U$$�3=S�q\$|��I��R-�R�0y�2H�!(C�򩗟bҹ:�����A#����+RMA�\�˦
�*N?�Y��,���O�y�m��;��jF�����e��I��h�*j�g�FV!����y���42a��P�15�hXH�¨�ݝ��K@<�]L:��Y����:�� (Z���#'}{��W�"0�7��*�2=��w�FK��J���#{�j�"[گY�����Z�O�Y��ܟ�(��lW���U3� a]W�٘����G��/1-(�_��]J��I�l���7�����5�s�J��[쏤�Ҟ��.�`���M��I��s�	˃5m���ι�K��"��M�Dk�������R�FSi��	x8�E嶍2W�q�j֊�M���D�T#F����Z`�X~z-�훢~;�@.�QU��阵���(hy�F|ᇩd]3L��y�b���������R�XB�Ԭ��%	H�Ԃ�6W�B2*�6�ذ�$F蕃�>~x��p��ą��
3K���w��p~���2��&�-n�h]�$^��$����{y��E�,㗁#6Zu����︩�C�P@��=M�[ZD �s}�U&j~�ă��s۟	\~���B#;�X�3��zNb�R��ӑ�0�+!f�xw���'��mP���W�Ҏ���0Xj�����K����\�T��W���������|g�V}o|��b����N8f�BQ�'���O�U,=�U�ŌOe���g�eBI]�U�~'�/tH<�5C=ۭrnށ�V.��ɧ�V��G�k,W�+���^Dr��4ʯv��ͳ	�X:
5��8Y��^��,�G
�!!,���)`S�e�йJ8>�AX;u��3�q�<��2al�7C2����ȯZz��~�~	Q4ʷ���u�Fu8pA�&�S�"!�V�o�B?D<�ȟ�?�K�z�����x�#��5TJ�;3\�����
�e�����j���{���@����#��B��^IHh��5��5����|c�'L���:��e�'���5�7d�%i����f�n�;�f��b;_�F2�uͱ;�"��4�5*��)�/���Cw+�9c���ߦ�*>\���@\^�VQ������A�F(��ܻ�S�s^&qi)�BЋ��	��#Z0�m�����h�,�#8[G���|�����.H�O̐Z����[�ڟ8���<a��N�Vl���+��!+�P^����i9Q�N퓔&�\��Ȟ�њU����)T�.[O�7�o�A��s�0Q�@�9��	b c
9��sPR���+8��K�w�{_FIo�y'?H�#S+�vv�{���N�3����:����*�l�q/z16�̇r�T��y��C$�Ua�p�����w��I�J;;y�B�:0�@lw��oveL��F尟"��)9x3�	U^J�eQm�h�8�G�V��.��ʤ��t��#��PLw��%>���ml�홅U�*C��/��A��0Vy���Qs��;���O��(�Q�Yv��
�*^*t��bL�9�#M�+p)��@��8�|؋%��Vq��xnFF��!��8V����ޑ��O\�W��kH����j�F�zk(��u?r���ڪ�wR�K�v"~	�>�"_-��Q]��$��7��t �ټ<�����"Uw�+Fȝ�^�v.h�쇜.%���y3�o��[�dt���G`r��_�=[�@��1���u_�A�e����<��30���>J��MDc�� p5%��ݮ���l�Bn"SO��S�?1��|�_O��}�ܜ��/�nZ>��4jS��ߙ����u9�P��f��(yܭ�`)�.(iYj2v�bH|�v`S|<p��x����9����w�zO�1�PfL�tv��/�J�όl�:L�Pu�݉���
�7���`���_���0��(mo�z)r��m��Ze�WWLVs�gp4�(Rx#��H�Cj h'W7��J����*�Z�͢�6���:	�=k�e�.[<L;d�#�b��gDs$"�A��G����x����.ʸ�T	��h�Ŝ�!3!*�bջ���E:�xa�ZjǴ3�O�7�2����it���~�,�g���"��O3��Uay�����dı�b#�wl��2��B����8�*�u*BGck�S:���q#`� @O�6�v<�U�����-�)@�b�襰�;
�l�d+.���<.�=�hKw��c��p0�ul�f8	@��i{��SY�ŁG)]ٟ�Z���i��P� 	��[.v��\.�/�R���4	�̨���_��%1�5�8l�����ԇ8��Em��vd��gT#R���NP��:6�=2�vXj�F|��������w]��eI�ۓ����>���''�
�� ���v����l�q���X���`N�c)n:�ӑ����8�FX	��ek~VV����T��Q���u�mq����r�Ԭ8@m^��^�� �]�� �q��O�[qfږ1��e:��q��5+�c��m+�x�Ѹ�"r1���<W�,��K(n���~�q�,&Ύc��P�rOO&�`^���g��MKh����t�����<a���������Z!�e��_��㧓�|��2[�Ϭ�Oނ��Ġ pK.쀖v�^U�(�p�~i��<��5�C.y�~��8���T�VcG��.ٞ�t�;C�����?�í>��yg�vff2��1))tC!BW������Ψ��c���N�����\g�Z��� 7�Pc 9��Hn+�e6Y�R') ��5�(P���:[8�r����r��H_��;�Ǜ�*��:�$�a��+z"$���kdRy� ���e��'�o7�>��a��5�#�q��H�4¯��}�9P�K
fO?���m)Ϻ+�n)R�5է���Q�N�h�;񲷬cybww
OrY\�i�,��m��pkx8b�ı"0l�[�G� ��]�����!��k�?����g���ޠ 1^�����!��4Y~��A�e�ߒ	,�*;�#�� �\�fM�&]�������o���45z����?���yi#��.���4��u�G�4^pbfuI��w��t�a H�UIGk��(��:��3Z+Y�j��
�q�d Z�Oz�[��+;(J�g� �z�Wo�j��5��H�q�wux�ޛ`�;F˷