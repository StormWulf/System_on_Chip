XlxV64EB    54b4    1000�����h;��+t�a�mT�ݰ�3���ul�Z����ҋ�/�x>�>��-�� �(�CA�Up��b�+{�óB���(z������0�������ry�n}��Z�A[\��=��b��o&"ʙ۷�lu^f��S�,�4ܨ��h�b'���r�4�\�=�J�oв���M���$�U���3v���S�nB`�X��I�P�������H���cߏ�&Y��O_�R@ ��j��Շ��u"��5����!�Q9<� )g���J�:��Q<�vD�t�s�h��YwȨgy�� ;��>�O����4�SJ_�	��l�iu�
0â[��L�7��A�u�fc(IOM�z��	df�N��bTEC=C��WEY���+0�׮y��v�Ob$�@a����"?w�-���|4�1�bP���k���%C�L9��d�;p>U�I�H�'���������1�&��%eH~��o7`G����]r��DV�A2�a
� ��<��{?�ɋ���F��*�/񚅝��"DQJ��w�>�\�JW���e��q'�b�&�g}Ih���hI����H�,���K�\�{V�Xz
�����BS�=�+���:�������\CL��B���z��Ѐ:���M���B�%��͊��f��Td��&��̯��@����nD	�Y)9�%�����Ԫ]����V��f����>����}����R�2��_�GT!��8�՝� hA��0�x�w ��x���-��#���p\mt_Ȇ�K v����3�Z\N��*K���C����ӵkJ}���:L��N���/�j!M֞���"kmR�ɬx�8/�!>B?�� ��LK�zmm�Y�l���E��]IK�wx` ���)��8�=���	�7t�� I���b���ؘ/��P�D@�E��Jx�@"g�У�B}�H'6-s[+�
����.c6%?J�*𺍋4�9���ѹ��}�f�:��V[HRn�+}}�U1GQ�U,ܜ�+.�*�&��/T��`���-���.K̞8NF����/��M@Q�������g�?�L�� Q1J�s�'�B���p!�U�с�o,uy%k|�˾#Y�c���uG7d���z���|��&�X�B��wdĆy9/乊�5w3eT��rk�5MV3ѽ���	n��ü�� �K����W@����Vr]ϖ��{�m߹�M%#7�g<<���y� ���:����D�p"�m"Y��_�b@mut!�.���T��\�V�Ir��#��z�%. ��<��-@(��V2Z>1qB�+��a��$����Y�<���k���8�I��i�f^��~��迩�wT�2h�?s=���,<�IԔ�~T��+��/�dS���BIX-u�r꼆R�~��!��,cn�$�fx���k�Ga�� ��n�YT�F���f��~��Yl�a�$����`S��'��DP�~��߾�	H�g�*h�
�S$o�~4�ܸ�gw6�v)�8�z�Y��fG���	�D�	g�&⠡�]	�[��&��h)`�\�b[�Ӫ��|���|j���k�M�Qf=�$��X�	�2zM�@��F��|]���d��-�#�D`S�f�X���ٜ�tk��s��P~�|��8��Az�A#�#���#�i��B6"� Êr�9�⫨VB~6/6e��K]绥�#�ĥ}Qq'o܄R<��7��LV��2(��fs�S�j��������,������mЅ����K`ZV�O�rL� �W��4dK���*E��+ۇ�On�8��J�ӓ�X,/�ͣ(R�-��'����ܖ%}�F�L��`�r��fک�w����)�V���u�m�P��`���d��)EU�;9�&<�Ѳ!X�cv��d\�Ԧҭ��	��w��[���*bS]�(|�����C��W*��?��,��?�ܽ�.�p"��cI�j����`�.
�s�V1+��ӿvC���b���N���_����muX�;b��Dǆ*Z����"�#�C�S�ި��D�_u�?9�JU2���e���Y+&����}x��N%�_�`��v����|�S+BY���^�7&�m��'��(B{57{�
�����7�Y���ݸye�֯\E��}f�j;8V6����e�^}�#����Z짯��(n�vqXӖ^t=L�	�MC�E�dNIÃ��|u !տ���<?��0�L膵���n��I4�F!�����bGR**Hˊ�
`���|�B������!z���*�=�:!�~�rq?U�A�܀��r��T!&>!-q�-��z�/��^������2� �@t�r͚�����ԍX�����w$l���X�ޙŜFb�(?<��1�k�-v��\
ݚt��}��&FO�WaOFv_U�nL�ڤiy�Z�D��*j�u�� 4n��|�s:A��,=D��Ӂ0��C����p ��M�̊����}�6�`:<���U�5;�`�A�W]��J/�u�IKVJC�-G2Y�珓�fI�/��=
����a^���&�쇕�#�ל��+T�o���v藩	���]C��$^��tohgo���W"����2{���>v��"������~����L�J��b�)b��Q �\`s�+)c�T�6q+`���~a�桡&oˍ�"�,v���R�R!f3���ʭ��ګʽ�3����j���ueK�S_���nK7�B��2ϥ��"!�U�Rg��!�%�:��O;��%��l� u:��Ѧ���j�Z0���١+��і�G(�����^���N��,R6�E��)�ߗ���'�^�f���3ۮ����v��S�[.v�3Ak�����.n�P����ǫ�I�h0�������h$��M�����'\σVF�M�'H��B���*p-�$�z��Ш�"JŦ��4h��ݸ���If�H͝���Z�呣�Y�D�ro����A�zZJ�J�I6��B��TR��2�WU2����
v�֊c[$P J��#�����z񿻮�\�4M���r&�]�>?��{��ͮ&�Z�'��!�����u�Ǻ
�ڨ����v�ɑ�D��3�+�9⌃��=F�jz)�`O�D�Z�g%�H{?^%���|R=�O�F��JX��ƏN@�@�\�.�f`���P()a׫���d/���#�`�ڀ)��ݹ���nh�����>�sC:1:����J����C�;�{�����c��Or�Ns�BN�eJ2	�Rv,&[ �\T�f�z�*�O��8J��6-������h��A�XY��3bE�p�A����DV	���nK ?n�S���ݥu�`ܡ�?��Ϡ�[�����s�@���-2*�K�Tt'1��w���]O��6qS"��)P.A�rXߣ�������.���d���q����1�")\j}��$A4𾍎N��ْ�k%9�4at��y�r�d���}�L k���"hl}g��r����8����'�>�DL9+m���#�M6����2&=~�� ��G,%e౜��@)e}oٗy�ex����SP'n �	n����:�%%����HbNƂ.�~�eH��ڷ���y}1(��P���#��~^"�:c� ����c5�0iDaH�@��ҁ(xX�M:�@O��R�.���Z9���m�a>���?�"T�Ȍn�T�ץeOL�
�5��Fav�F�iB�>A��
��-��R�"���]�n����t�(�}��h�3�Z��"�RK؞ �8���0z��#��C:k �<��V�L���Z�ԫV.�?��I��$]���{�}hY�ME�w=�l����P,+�Ӂ-���&sC�e�ɧ7�3�w�˒�$q��j��Nc��B�1�������v[�GB3;�^W�`�T�Qn�/�/����rTL<��9�!��kYMr��Lc���G�ݚ��%��7ݩJ>C�4殾|(ƺ���e�w�H�V�Y�4�0�P;�"3w.! }̒b�R5�a��z����l�@� v}�d����2$���'