XlxV64EB    578f    14c0� <r���Nɔ������
�An���:Z�P���&�ϗ�E|J�o�!�̈́�~�hwI6{��|؉"g��|�)f��s
���MC\,"�"s�z&"n����,�+(���w�}���!ɳ�G2U`� �a��!����F[B���R{'�	��@������(�F�G���f�Tc��p�H�T���o�<�jN�2}��0��������xI+���� �Y�.��)�t�M���q\�yz��>F�E-F�i˷�|W��o5�'������v�e��:l(��x�	��S2t	���t��R,Kٰ�qmx�qW�ܒV��I\֍�V�����}����z��E�҂�� 0w���`����ǥ���׬�*d�}/�X١M��iVL��*�̢�ˬ������[x�:�Po�ry-"@�!Ҟ2a�A�ԅ���=0��z֍�h%�dR�0�h%��N@l8�dC� F%^��#_�������C";]�ۈ�q/V�w��I�t�(@�<GĶ���/Lt7�@y���k}LZ��D��P����΢�:$"�����9CP=�L�x3�u�k��U��ѥ��F��q�~}ݏe�C���.g-^p]��4a�<=]&)X	�,�b�+`��#*����d�)�Ch�����y0��,׵i̊��4Y�i���n.l�ն80&�D,?X�lJ�T^=.	�swQ"7�&MI�Sͅ[P+l�8�Ge��oAU�pUv�/$`A�$ 4�~�3/�Ny�i�Az[�mT2o2-߷�H%WC���x�����4Ө�n��~��gx-l~��}��޻4��4!��8��Z��yw0�+ &Q/|�_bu�RZ��{�9�|P����&6��Ӎ�9փ�̛ډ�&��G۹,��\TI��A��#l	�&�/���,]�i4/��b�/.ۘ}6����d���-�$���$O��?3A�C����!�zVܪ�z��T�N���oAD�h�آ��\�bi9�=$���$,ܯ5B��O���{(䆜�o�����A���i��]�=/ө�oL	}>[X��e��W#�F�Ժ��p+7�ۂ��uN^W0���Ȳ��7��Tgԉ_�.�Jwu2�b��Ax:�D9�
��C����`S�~�y�����o�|B�v�;�h��
��}���#���9 Y ��c#��x� �ا���*y^���{T-�xjF��y� ��(��E�Y���
��>nX�a�����Jhn�y��$��m�ꠋ��Z%� ������v`�[�K�5VD@���O��ٰ����d�z��t4�[[)�޳ğc�B�d��5��z��@=��}m)@C.F*3��<ǔYQ�,���s#�Հr��0zsߊ���+�](G�����+�ja�7���O��JE��+���)h`� �$;�#Qx�fƤYR�j)f4}�5k3.������\�[L�).�u�s�9	�I�\=�'j9��Ci�1�HXEg��Q݅����
��,ߧ�&L{�Q�ShmNa�������:δba��O�G�^f.SƊ$����!d�������`+d8{�8]��6ljwY�|��S`��<���si��M $2eN��\ل�y�BƘ��`jJs�I�N��Sd����Z�"EhO4��V��ߺ%�Ύ�ȕ|�!����$��~�Y�����R�,�GУUoQR�|����N{��MÃ�dBH7(4-�A_O��L��ۜ����z��(����Op�4O*(���c���|��؜,�}�啓��0%���8x�eq=����9m��܏o5䜄C����Wx.�٧�����<p�`���0�0^��fch$�ٗ��\	O<�#{��g� ��t?����ƾ�aO���ƕ�s��v
�{�7r���!�6ncI�kDKP�c;F���qק���l9��ew��|_��j�v�3��Ϟ�c�f�������N�V���}����]���؊CD�!��*�r+��u�]�|�~�x`�f��|H� �5eK}L\;Y?��i�~�����]H%�P�	2Ƃ/�l �:�����Iy�/8�d�舴���]ݍK�m��ta�̈�A��f�1��{��2�}��Q�d�ƀ�򊍜ߨa���~\�=-�3��4�_���^�s�ϸ����<$�ւ@�M*��6}����L��̛Qs����jSѨG�VP�|`���0��Ⱥ�I�k<#�+�J*��n���{OV>>�	o��ۥݎ_=f^��{\�a�?C���SIy�� ^=P�-�{f<�D��)�U]�R�$�@l��70�:<��`���%\��J2��K.�a0:	q�w�̆!����a��r��Μ�6	��և�q��&�qGR�:d�G �룘e���yu*O5����vx���r� ��R�tl�����:t��'/ϙ�p����6�D�Sv��ٳ�gf;�Q�k��̧�g8:���O�2�e�˂��
���~[m9���/��
\e�ۚE�B�۬�_(�����?p-X������)�Wr�T%�̸]��b�7��	e��$\d�W���=#zsK.T��q��|3;��8<�>��������wp��`]^-��lq<,��wq9�]h��k�tC��L�Q�M�|��Չ�i2���4c��Q�S�I�y����3�2�Ն�N����2�.	'I8Wt�<d�ƴ
��kX,��t�*���<�7<�$���ۍ�l8x�CD'-�G�K�]G-��.���E*Ǡ��ʔ#�wA$�U.�_���(�ٗ8��m�4�����b��F��EY}�ًN�Ʒg���v&�wb�����=���5,��S�$����_��j?efr�3LJ3�s��Ǵo����K^.*q�p,����ʔ�=?M�>��oƝHQ�:ζh�����1-� ��:B���;�p�_y���)@�{�u��e[�����B�R�u��}��J`��o#hH׹�fj��T���%Ϧ¤!ӂXv� X ���,F��u �����!��k-dd9e%K��BM���P���r�O�}�tKSμ�*ߢZb3����f)Y?C�VnW� ������4;���N�D�ݱXAܠlV�`R����C�Dg�|�Ҏ�z�vp��6lg��y[=����>�+C�
[dE�3@̉.=8L�ੋ�C;����',-��b�q�C5Zn�~j룠���7>t�����mBф�ǲ��$t(�JEQ�ӑwH$�p�{/����f�bNp� ?L�D�T8�N޶�:@�t����e\����4)�-�T͚�k�H 6/ ��etAɶ��"�?% q��QV��É�J�����sY������'zi	��ř����$-U^oYH�r��@��,�pkx�S�=\/+!(3z�%9�k^baK�t���p KIױ���ମ5r�(��K���5T%���7�aw]�[[@��� �"HO��#8dwԢh�	I��^CG�"���>Q(�vzfw޹5�̛����F ����K�[ӱg�����IM~�������OfJ�]�l�a�X��WC$%�Jn1f�B&�,*���Y4���|�ˣ.'��R%zA�v_b*Ӟ���w�~Γ!���8�lN��V��S�v(�Qm����?R�0f�3�`�M$P��lL�^4#e1/���C��8I�B͜����y�K�x�6y�><���V�s!%���@��vӉ�R.�6�[T�f��bi���a�?�ɝ �a�����26�����W·WK]�ܠ00q�_x(1�3�IT���g%�BOg	#�qQ�_4]f�n���^�X�wr�&��5���}T1iwP��M�i�W̼�n���a�jb�&He��w+���P���~����M'�$񎽁;���OM-�s1|�=G��dsYіo�k���x�� @[
�<��.̧\ByA@U9�d613!��~+s�_g|̏�܅O� \�y�0�c��hzr�+��H|�VU�z��,%�'��@����*��d6пL����������ҕ�j��|��b�Z���*��W�f�Y���_��1��I��;��T�p�oFX�NXT
A���ly��PH�L7ƭ�a僧?		�l�"���!�� �p��O}i��	�3Oqf�#���9B��SE�Z�b�IT�������1^��ĭ�����,�Ч�-����5�R�T���Ḏ��u�i;Ű�A���H�6�iIdB�pYv���J�uJ*�>�=���A�U0�ݥK�����CA�Ӛ3��2:��Q���G2��w��샶�/�a�Z�*�Ƭ�)3�VȄ�{���((��9���|��apF=U�e�Y�X�!p�9�G����y�	O�N����Kz��A&#���eV�1|LB��s�5k�$l0N?5%�O"��*0b�#	�錦�aD;)>�ß_�B�{.�CV��!�e���j��2�R������}��l��F����D7���!-ĳ2"}�lJ��)�L�k[��Ͻ�6M�=��eq9(͡���8P�Ť;��
B��W>�o �a��I���`o�iH�y�o[�o�9���i{�����8?K�6@k'�S߻vE�a��|�#��!�Bg(8��2Y���80n'8\@��\o��ߜp�O��vR�F�5Z��B��V����F.�p3������QKԅ���ĥu�g#Ղ���"�D��K،>
�ut���H���CP&u���
��o��2��A�v����.-��33����s�w �f\2�-�)ϗBo�إd�ᝠ��du����3/��-M�m�;����9l�
L]����i��()<�G�N����AT¤��﮿�PZ*P�'�l�>�3�"Uu��C:��o=c����Z���p �Ie8i$u���c`ٶ�8���'R��]��v�]�&�RYX��u�*�%�Ha[��WA�����+] �2�O,%�b��"�3 ʡ��L��`�|~�3")���:(4���%��U���Ǣ,���^� �[��=v��>ZS����o�ڤ~;٤�*pJ��4�?'֭d�#�/���Y/�$��M���X��Ń�l�V��Cӏ?X��I��$��(\�
�X#;�{F�v:�j��4w��j����T���/���~)���ҸG��V?w�4�D �N b���~