XlxV64EB    1f60     9d0�rK?���8AM��9�xҙ�YV��c&�r>� �r�jH@	����j"�K+P����vC�L�D�^V-�H��FÓ��F��'��� �L\�V�{���*�\�X���DO��˼�u�B���g��4ET��q��ѱ���Z���>�
WMG�W���K�^D����*�j�EQ����,�J3��Nf���x��i���"f��? y��B�-'#�%�$���ؗ�C��~��{�.���Ns��{;Ǵ�X���C���LB�9�������M�ULh�]c�f���B)�\�ۻ/<���W���fwשZ��Ӂ�8��.����E���	��g�u��)\U�%�A��諱�h���V�dg��O
��-i�V�F�h/��d�VjR�
�&��f��i��~ˮ~B�X|V��-����4*�]��d��#j�5ֳ�%$RuYn���=e� %p�'�S�����6R��h�P�ے���;ñ�D���kwĭ���@���z� e�0�����O��0���|��	,��0���������q����9b%�\G�˄D��i�_�Q̋ޗ�=�Y0�.2��E��6�~<�k�xW����H|Pg�o{����	�:*�S�L|�Z�����FR	7���e88�Hp���9�������\c<^�V�T�r�管�b��7*�R�)����3Z�4�s��#���}~�Yl׫���_f�
����!�*uP���ۜ���=�_�5]�
��yA�7v���R�bP9��~�~���#�,��F�����͋@E�;x��)&����(��'!b�����a
UM�-� �!����c��$��[Rmv@��1c�
 �����*]<hFI��[%
���w��D�_g����6��tZ�ǌ�p�e:u,�<�#�o��Q�Ė��!n���а/��*I�'̈́h��w%�L�鎸�F]�� 0���Q��˕���WjL�J���v��S`.���,,]�R��@e�$�������"�i�*�R�w�=e��U�;�h+�%B{A�oҹnS�<�} A6S�*��W�Td[t��6Pk���b�qQ*��}��e���C_KSJW��nځyx�������|'C����ᐜ"(�'1�� B��ՙr^6�?��mR8~Y�$#����,�q�~����"RC��[G*˧k��dAX��n�˧����b�c��h��6W� ������+x$�1>����EU��О�m�� *鿅(L{�=��%��|W��t��ҟ ��ɩ5;E<�9y���[�N�SǞ	�ŰJ/�R����M�M�
h��٪؀�°�aɗF����<�,ȶ)�m���>AGwGG������v�g9-\H�����(P\д���d��э G�-|�)_�F�b��F0G6	h �Ca��跘Pt>�ه��w�{�k{�dj���h��U�<�^j�c)��),D��7��
����x��5�V�jN�v��=����s��B��0�-ս�2�˭9d�m&�G/��M�sU-���S��V�3чQ��B�(���4$@�5[u�Fyf�ĲL&��>D�F�uw�����H��f
qt0��N�(����1�K�1nBpl53{�ê,��T���*X=
���]\<u���ɶ?K�����"��5c+�^)���X��vcN��k�2$7�A�yr����:��o������r�Z�%�޹=vP�I�#�=?
�"/���8$	��s�&*�q��]6� jh��S��	y.�?)��dG�b��W���tuQJ�y�z���cIF(�_7h.KB&�HQ{*�[�1�O�rZÁ'�j'���b#a �pHΎ�j3e�������W޶��sΉ��+�+��R��𱓺���xBG|vE�������I�9>�U
�!���m����q���B��|F��Hkn�.eG���F�Z0��?����e�8eT�᨜�ձ���j�����G\g�����R���`}&-ńc������m�4 ��-[��6��U��f������X�"�A���B��IM�gg�,!}G|���[z�|��<���:h�z�Y�����O���>��i�x�e�2���
���d3������%���,�Ø\/S�r 3x� ����e32@?~����=��-Q��I# 9Z���!'J^(-��S�w7{�NS��
�ʵ�o��Z\�5�F�����h�u��Q�6��욒� g[�{��y�h��:�������=+-�d��aH%��]f��a��룸a��#�z:o����杰�__�8��/9��q�DI�?Z��Z?��^O)C=^��UH�c*�!Mf�F�1㥀]nL��gr��
��7��&��Q���4��)�+��t�����HjI~��в�:|�s#���l�����G@E�ۮ bC���=Y�o����G�%̎�(����G�1pkCE-