XlxV64EB    18ce     8f0Y�(y?��H�A�ta��aK�l���=W5�=$_�V2\�bb�w�,ܻc�D9x��&�}�j�Ӳ���ƞ�j'���]�S�kE�,7h�Bt�`�}����דS����VM��a�)GP/`2(lt��խ�߫o
=��Os�ӌ�T����BEr�a�Fv�����s����b"��H�Ӓ"���A
�s��"/�U"�B�[�A�=/�m���!݄���c���kI߫.B�(#���znI�"�hܜ�5�(g5���Pe-�T��vs�iTW;���.��)� [����˾1�a
_X�v�����R!&�=K:��`��5l������?��[`�x��ز��rֵ��oW	���4���mz`�>Z*:T?{x����A��s��	��/�GD��[�\�b��� �,��D�'ʭ����q'�ѿ�T�����	ƍI "��"9ă� 5�?"gB�k���A�w1�Zs��$��\�Yr��B���5|O��l��C]���B�������7��~�z�K�U����?�+���K)eJ܆��v�i�)s�1	��L����I�3`d�/��G�������.&��2��t�I�Vg�t"�_�dlTfۺ������ޭ�\ٸY���^R�H�7�K��ֵ��h��|�������'�!�(��F��EƠ�O�U�G�G@�����/�pr�Nz��2J|X"_K��I�v㠔���K���K�]�"?y����'[M���!U퓙f�f�c|���@�m`��J2!ͩ����V��]n���s{zL���[#ܙdT�w�0k;r��r))�ڻ�MU�9�~h]�I,�,�?�'�Vv�I���|��0U�W:#�UB:~Ag�F���t,�.��2;Ww���^U�`�wΏ�wb�$x!�T�ѽ����s����CJ3��&/ε1�i��gT��C��0�yzq5	�_�d\5��Б0��V��z�5Ҷ��]5����f�t��3{u_&������թ�Y����'UX=;<�p�[�)p���8�s���a4��LO/�6��C����5��y׌��M�H�@��j�K>>a���F���8��S�v���K\���ZQ�q����R�3`ހ��k]�{7��Ȣ�Q�Z>��*�W��m���Z���#A���=p
2�)����P�������YB4��a�GP�t���A��f��5�@)�cM�]yZ�	9�.8�j���7z9�����0eos�g%T�V&�6E��Y��Ӏ @;(�w���M�-��?Q���:ɍi�ͷ��D������t�#D\ ��ux���W�&��6��nM�	��q%��,�jZ��P����>~�m�p���q��������56�����k�|�ޓ�����(s���W�Vy~� P��:S�w\�W�s�θ*o;�z�nD���`��@���9�|��z�K����"���šf���u6AcRD���4��x_xn�yqpp��J���!,�BiA7y�79�u��췁�i�� �p�h���C{�K���U����;<n�r)��,�z��ތ�G����$i@+ 3�G��e����(�F��j\�	1�TwD|��8�ed��(._�Om��I~��i�6���vDQ�A�	Ɇ٥�XH�T��T1ɬ�W�lڧ��5�Xg�U	�P�`W����`�A����хmǅf�z�hé����?G蚮������m�����zZ���I���Ma_�R�Ua%ݨ���G�_���yg|)�^&�r�#a)��-L= ������q�d�a&ۗWY���L��������ώO;���E	3� g�g��z��BS�7���Ex�\M��V������®`����d��Ƃʣ�;vxm��I�g�mi=�"�(��
���@yJ�$i#���w����̦Sg�K:u�R�T�����agW���l�*Ћ�$���������vwmz�(��.D��( A�94�B��ۿ������e�m9��J[D�*���v�&�U1�B�W��F�������U�n�kC��Fu�F*�pEbRi�$d��>�8�PbS,c��{C����h�(Dƾ��h�z���e�A9��2��٢���6/�O�
g=�'�ɳ��������_��0N, 6������`��/w�P���F��'J�j��`k�E"^`a�Y>���#|P��-��<���K~rQD|H�ω�!��I\����uY�k�� ��EhN8.�U�AW���