XlxV64EB    17f2     9a0��/�4�&�|�ы�6#P��(�����1�j_��U���w��dV����sS_�a��B��B��$D�]zC����ױU�ݭ2=_G(UW1we��s�9Q��G�{ΤA<��Տ߫S�&���s������%Ԋ�{҆����9(�i�;�GQ�rQ�������CO�Q�S�Y����5��$��4wr�6M�My�a]7D��Y���?gZ2��vc��d		v'��h��֭�6�Ҫ��[�8b0�v������.���7ZCK���o�EU�/�!�m������q^�5���ˑ�,ɇ��c�����=��'0ʕ���ȫo;u��r>�8���&��_!G�N��/N�2QӐ	BRR��a��Cت@�?��j��Y��� ����m[aC>d;��v�_EYAV#E&��&+3W�B=�C�	�Ā4��g(���{+w�����v:�ߗ¤`�\t@(��6)�meIݭ=�s�)Sr|,MMkl� ��D�& ����9�M%�'R�wqK�tn�@��GU1p��q
���FU zمKy�"�]�m��zň�����?v�ƞ]�`�x�Л ^�mr�	+��ЌZM��0B�t2�~��	1����$�r����q�dG9��WW�k˔F�o`���U�06��5�Pz�Bx�X�mý���KB�(4�6X���T۠| G� ���e���Y��9�'�����ڢN�W!�V��Yc�o.�O�z�"���ܡbyޫ��'�n_��q��MX��=���|+�ä��H�^C��G�a�JФ*+֮Q8�L�_:f�Ǉ�~�� $��]c��v����q�]�H�]>��S��~_HӰ��i25�K�%�޹LJʤ�|����]���藾�1����/	�j)XU�d�'O�!��On�_DH���Ά�5�|�F �px�����i�5<���cS����*�/uh��K_��� �
�ZrO�y�b���gHN�Z�Y~m�ު@��E�j�3a,�������Qe�`�� �ঔ�G�5w�qbdyg6������,>��%��*-BM���ue�
�l�2��U�'���w��V�k'Sa���7_�a��6o~'(��f�����(��#���'[��U©4��ĖG �]@<�۵CG[0n��/����󚤪��2�ֈ��oC?��MF*\m̢�*S��>�B����e�yvϕz�UcXН�S�!�x'o��|:���%؆͊I��-���Gh�����p<$!�PM�l��ߧ6Ň���|����[��^C�o���
O��1g?=�'�!��j?��������=���!�Kr� �m��6r'0����pA�
�L�����ԧ��kRC�t�ȸ8��w+�Ynm�H2��>[IMl,�_�n���� �-���*F���,'��w�o�g��0+jZ�V�)'�EC�������`��m]��*ž�nj~u�v��S���o2����]>�z��E<� ���[8U��+�-��6�n:׏�·Q
E����� $�v�X��}��*ި���
#��,@$����^�~����N�����-(k���3+hr��Պ^�z�W���,'H�^�x�hX@�c
*T������m	�Fqѵ�,U��J�0mñ�s�_@\�:y� ��=v3�s ��*&X�Y���gLq�?��Xt��g�)�Y.�t�e�0=ȳ��:�Ҵ
7��g�}�H�g�U�n���ꃏ-3�ަ���-��B@��3��%����D�C�]>ksn��R�"~�	�GE ��j�sH/��Tm)�-!RZ���X�1(����;����R�I��[�$nſ�.=�X���X�~���=�-��1�7�wX��U�Ж��@~j��1#ܶ���8M�j��k�Y���ec�%vt�A��;�#{f�cV�z�o���|������<���-�÷�z
�Ԝ��f	�	ĔLJ5n��-$�����m;�9
�gQ�dMǖ�u���$���ꗖ�9�V�����ŬA�ǟ�ܵ��]�o�����;�ՙZ�A��t��H��J���_����n˪�� ��xC �:�LH�CY(Gi���A�F}�}�m���"��H�i�����B����ƵS�3�혬xk"[=�|�E.���=6;��(�Q��j�xicl��:���]�����W�ԾCc��[�:��Q�0:OE���Z�
"���J�|~p9�?���	Q0��~��P����_�|�d�MU� �7�_A�/U��5�K6��y\*lA1�Ub�"�;�L��� ؊QO�B����i�G��W⭌�à�hq��C)�������3 �$����b������F��
(���l*�a�����{j3�{.�/fy�e &�k��d��k�E\z�6;���hy6S�b��F�9$�qd�kK�������M�;4��h�{�]��W�2���$�FG6ZH��Ø���y�