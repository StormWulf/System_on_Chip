XlxV64EB    fa00    3010�^�`[)��[Z��VU�9����i>uAD��wQ�2�X|2o�'��5%ɦ]*t�׼X�p�yn�j��n����(ߓ;����qzpC�ė��ǔa�#km�+<7�p"�P��sP�oҼ��錀�Q��}.���!r7��GI!t��zv�����9h�Gy�
��/=���;r�����[TB?,=u�:�+{����X�EU�d��Yurf����������{IG|kF9�]t)�{�Erd{z�wР����^g5}:l6���mݣ��dA�{��>�:�p�+XMF��il�qʰ��d�� r�Ɖ���nvI,�x{�������dɇ�P�� I����GD�G[��0���B˳
W�pU�e ���d!��k��T&����X��͓���,��Zo+# P[	4Y�e��v�t"f����)&���6�a��ɯ�b��~AmL;�����W�-�[{��L����1��9�����eŎ	�[B��V���q�aM"���ig#�h5��0�
�.�[Xg))R�}����׳z����=���r��0�/Z~˶�
�k;��ƫc�]Oj_R0E�4�َ0���
V��H�:@�����������a�����;�ġz#�>b@������H�؊5s
9�ؽ���+�ާ�]ب7}bz�_���� M�<�ɣ��sD`�:���:|�i ���Җ�6�{���!�>��o���Bf�1&����a;&rk�k[�|�7řp��4���I�~)h������^c��uYZ�ث.w�0@� l�r2��6�	��o�����gڽ�3Wѝl�+}�z�x"���%���sx!��ɅTφC-9VC��F5�2�o�H�������D=q��0�_�y��Z�͗EfDK�'������w���Vݼ؟��=�a\ψ� ���٪��N��� ���Vq�%b�a�5b�ⴂ�O�.��;0U�g�tS��V��TW0B�5���f��j��DW_��|?�HE�C�M)ү
�
��tFz� �����)��<4P�4�0��ε�H��"��0V�� ��]V�oV�'�q��;�/R;<����Y�Qb	��xy.1������j�h����8� +�D$����T��k+%Z��ђ������fߝ�,t''Ɲ�<$?=�Y��f ?�v������Pكvt!���I����6��A��0����۽��k�-F]�ѣ����V�����/�M^Xfn�:�h���j�jo���3#�R���%lAG��W�{�o�[�k4q��?��W��e`O��ىz��D�{����v!�RxB�#L�QX�e������iV�_:J�(H����1A���gR����Z$�s/��%��:t�d��X>2Ǆ^�/Es0�6�c��Uуݾ���U��^U�K�^��PR�����
�~k�(��@��*�eu�Z�
���)�Lv�O+�B�m��jj�`�K��2��^LAHJRv�~��4J�Ћ�;�a�b��D1Gq-��*�÷�m��C\��^�`c�t}�в��B^ bEQ�}O��M��+b� <!�0L�.f�@~\�q�EL2���8�!Q�p~��>�(�$8ŧBZ�C��}��0�E���N��Mؓϲ�X�l.Yǖ��RG�����'�z��Գ_Zi�RA	VL0��č>D��N��'�n����_�&�̅`1T�5ם�Z�Z�	y�ޥG�Q�GiJ�)D��]�t�7��2X���u X�2�j�n7G����S��"~��J���t�b���MjT?\�%7-bjѳ� ��pI�D�'�C��"��$��-����y1��K0�pPâ�	h�ރ�'��G)}�A���3
�n�ir�_���Z���=	�E�\PW����ȣ>� �'���0K�oO��¹6�j�)��r'˲A���2����WƉzˆ>d[�ueV9��'���";��Xd�'�c�>��]���F	����=���͏1���+�Pq%��]� �^������p=]%�;]b��#�QK����n�_!_�H)��?���m>�]&υ~�l��:`����@ZC�f��*s���k�'�t����{+)��|xa��*��"��,���OL�J��O{�<�JY�7�]�.C��~(a�7�y����?)4"LL6'���"�#4�>�vB����-*NJ\!,�i7`/���d��^'��;��l���
F5�94۳Qo>�� ��e=�b�;��V��lq{.{�����m������C�W<K��W�}�l~�'�R�0�[k^Z�ZcȢ������ɵ�pN���P�������x��ӈcT���_�	��t����H%��o�6�Э��"�IL]cg=d��b6�{7U�9L�{��n� �_b�s`�Fct�/��r;�3qL%��/���G�X�
�~���(��'~[�f�����*�H�G$J�R`�V_�$t�6JG��0�7�j��)�M�#�����bd�&��C�a�F���6�Y���М�1�o|M�hr�n��#F7�x�	�s��`��M+],=�X{�ݺ���1��j�ކL0Q5l�Wo}~H3|�����6��nz-h�G�I# {i޾ղ9���H�&zNy�w��0���ió��Ajȷ-����K��Ly���:x�S�^O�P,υ��>��&}G��6zgo�H ճl��]��sɮ1����c$? |�����M��1�(Z��Gt)�q��s�בQ�Ó?��((Y��ؙ�̊���9��_�E���N���GB�NEY�c)��G�#��]\R�����u]���*���S1� 4��95��2�2~m���sJ�<:�*��L��'­�H��Hb��*k�TFm�Xs���B=>v��N,Ɉ	��#6�S7��Q�ഡ�$���� XuC�5Gc)���BI�Yʙ�+��7Y����!}�"d 6b�m�==J���R` �XĞ0�!كg��56�hpM�R�����(�"�dM�g
fҳ�ª�O�4=<�].!G��}$b=J���t���c)(�ٺ��~��.��ĎB�$�,�p�}����C�ÿ�D���5�1�j$���IsR�p�zs��-�pK�!��E��!��F1�����q T�� М��b�^�n#���Bт��0�,�a�ʼ)�1��!��}Zc�Yu,����k���>�7Z��B-̄#��4A���b�����Qc������[���c���n/ă¤?ٱ����ǖ������WW������G�h�?Wsto�r��kR���*���lGM��l�N7�Q�V�&�i�i������r��!3��|-i��Q{�J���Xje�	�*R��k�_�iQ�4։�%�#�:�vU� �_><l�_l"�7!��lO��,ASP�3��u� ���>���������%�=$��R���saB�J#�]���|141��`��	�P(p:A�rc�#pϢ_PV��2Jd��W:�V���.Y����XV'��}m�#L�ˈ�~��+0]�;�{����N�kiֺW����Z��F��v�	Ш](�NB��/߯���p���j'�YU!T!�");�jNMZ�>L.y����$�,�q�&T?�撿�]�OK�v��K�3v�k�S4MV����b�1�X���o6�H۽Wd͎ ��!R���Ek���AE��ڮ��ԁι�(������i��{?e�����%�'Eoct�7�k�N]x�e$������p��VPn�)Π�dlP������'�s'��S���}番"4`��)_��o�h`)%E��o^�S7ޟ��h\�
P�Iy�Od����2T�Y�?��]_U�[yY^�VsR�r°��(�I�A%�� ~T�vK�C)����a���#1�-� \��\�uV���8��ǥ�0��h'�H�ߐ)ꇥ��[��G�V�i��ރ5>N�A�m�Y�[�6t�����g�2����c�v�Ta��A�v�������d�FO�Fna����P_ #�m�?\�y�D6W����p��[]ZA�;�"K ������r����X7�=-!M�4E˪��'\��嬛 �}*Í�r����-	WS<Q�`��~ͬ�!]^o�v�G&�|�w�&�+�Fw��]l^*-�������eP1vc��.�e��B���!�M K��GsXg��\��ߣ����d�S��Da�4lp?n�$��+kj�++�ѩ�ѹs���G���W�L����M�):& �����O����XxK�)�\���p>.XD����+_��8�2��OB������p���<*����Dr��������u��%�q�U��~`8�[�mm���NLc������"պh,�H
�
����nS�vA��Z/C�[��x��)��Rro~v��ݿ��k���$�c�9���E�*�OڧH�.
!{2���Vk�[�n�#g�P�7�Q<8*�{dG����q�&�JG���mq6|��}S�;�m�]�1�C�t����^��O2�yQ�&�+�������W��*��,���H*���Xt�i@�3�^��{���[0���_���"��Y��Zd��\M��]��GJk)��W�3����x���Y�ٮ�%�#�:Ǥ2��!޴(��N,�C�e����6��+�5���q��4�l{-��G�{0��`= ���w�㳛��>_������0�
7Qb}B�F[o��s�ȝ��P$�r�4;�A��|�L��Y��*��o�D����]<���a��p���%�$�z��/�mPM�j5�R�'����;�x;���n5�꼿}�B�-��zo���6�7���ER�����)Ɓ1������x0��X���=���zm�5���+#�Tc�--1#w&�Q��+v�c������ҕq�~X����_M�q���� _�ҵr`h��K{֨OqK+�+U��>��rF_K)�?%��x��p1��ͭ����W�L4b�'����u;����㔫���f��oK=��_G�?��c�8�7��\LZ`�!���t����'��D���� �.F��zPD�@�f���V�%������>2���'qҬ�6�H���>o<��f���� ��+H�_=]�L,"��ޮ����V$�������xy�?�Y�o)T�ǥ2���$䰴eS s�N���)�h��{
q��'i��|�D���$�41g��)$B&.������x�<�ޟc���Pcj&��EG�dcG�Yt�J�C�����ӈ~4P�=lCb1��A��=�C �*���٪�!�H{L_�K�}�^uV_��"X���3�Y(P7|�]ۗ��XT��4Vh�*,�AS:�-�i�)���Ě�fL����3Y$��e�h�0H����
Zmy	��e?uxj�[<7�Rk{8܁�@�ύ, ��ϲ�TJ�܋.�YKҐ�/�\7\�\�I��eK8�_	0A%-�Fr����R�$��s��o�QgR�퉢EN՛u���	۷��[���rp2`�+���YT#���1s �#��L=�s V0q�2G�*�-a��]��&�������l>�3��v���&�4S�C�^�\u�i�A��N�F�i��J����-<�Ӹ��F�v��DIˇ���r���ug��kgą�m���h���t��C�yV��].�,��ʐ
��F�G�1��%���C�>/�M ���(��犊�]�K����:4}�
�E]�Ox�?{*�R˱B׬���0�`��&�r��S�:%���o�
#�
���Ǚ�鏭'�<���=7i�?� c��d��@ڬ�\;R��R������g�^�:��<�|5����eн����Y\�d�}x�7�[s� {!C�'/-�_�
0�L�ɌC�J�4&���ԸD��AV�X���Z6\Z�e=~�v�tE��A>bt$^���L=i�>��I�t4"n��7�/-�uv%A����%s׶�����H��* ��{@G��>��'�x�U��5f�(͟8G�ꨪ��
��ӠGh�m$��ٙ6�mhG��F��a&_j�m�e��]Y�{H� ^-!;����v��h�1�%�H�ha(t؀#�$WAʭ#	������ܣ\�D�s���&r�ĩ�J!��n���5���p��j ����J�x#7�kK�a
R���δz�pP���-��[�7`A�`7N����kI� /�NR�yB����Ƚ�tS��Y 	r2L1g�ڍ,=��w^�$���S#�'��S�����v����N+@JO��C�թh9˘�p���\S���a�	�������i�.7�#�:��"�\cR-}S}���G/O���R��/mn
�An��n�Q>�а�]���P��N��˂�E�5lG������W,e��J�)#-�ϏV�k���A���5	�c�PP3��~���l�HǼ^�;��^����{�BKec�{�+ɞ����G��=�%��92��LLKz�ɔ�	'zjT�bN��i@g
�
�*�#C�����>�)�og���"w�&����E8���9�B�/ZB�7�JCW� {"$d��_G�-q��1*��?���S_�r�����V��*rӛ�Dǃy�����lyy}���y+23�@]��®�熹���a���^��z~�x$��g��t�N	�k%�" �&M����t���%۫	��A�L��Wa�=˹ǚ2�n��&!���a�a#l��j@:�N�H�Y�ƭ�����@v dK��\�f�?i-�O>v�Ȁ�D?ݕ�Tf�������*��id��9� 8j���8�;Z'}��޲WE�[�P?"=t��T)q����z%
S�MV���L��M�`}hs`�\\��Y��"hA�4��kF�&�8�4Z��F�SH0
Q�<���4��M�>2�`i�K�Y�	C�f�[���*^_@���5i�o":ۓtU���Z�>V�~W�}�¦�?P����HM�⠚�� �]��nD�LeN͋1���N[�Q���&/(y�LU[B	w6��.�D�5LD:����!f�����;���=��LM�inoW�����1WU�&HW��SI6����\���(�R����曻��5;L9X��*��6�t�7DAct�jrEwN�A��V�B���x�;���%,�&���T�G8���ȉ�`/�SԐK�\��GH2Y��@���;y����#J��	�0�i(��'r΂w�xh�g� 9T��Ci?�yDݽ��I ��<$K���?s͞#��L����4+��[둜��	sy�_�a�d"@��d�o�x�"r�[�{8��� K�ο�N?��MZ��*��>cG�5�o�+�w18p�#.V����{%�y�,�J��_Iځ��(ip=����k���~?�,Չ�=��S�����1m��x�w���I}_8�e�v�+X$�ND���yzPk^�*+�Yˍ��d��35<Rmj��n�1�7����1��XZ�W�f;�uK-o�_����da!G��Æ�؟��as����z��Y]�9�~X�[E�l��a\�D��\F��(N����d�/3_�Ӑ������d��[a\{R'�̂]h�-������d�`�W.j˺��獓0*ߒ��5��f7��MP�ĵ���*=!����o��u�`��@���ʂp�+6*��7h�)���a-��*쨸�.+>s[H��z=l������sH�P�h��u��s����)_q��&WGn-���Ià%�!���*3
���I�V~$��z�=���P�^�p��k����w���|��7�%��=,k� 1)>��FgC'�� �y����AR��BF���?=z:�nՓ����l2!� �a�s�-��R��gS0�gz�(n�3wo�ni��v_-�c�e�Omɕ��v����C̃��?��4$	��P�̅4�*?��~p���m�i	��5�'�w�f�
��k֙��=#ܪV��ĤY������(��m�Ꮚ���2u�鬿�t������V��_| Y�m�)
��"����$�̙ڣntu��6|���5�S����O�}�S�	a��a�s���Q�	e0�=Qt�9��f������6��m=&�t0pq'���0��F��}�*
���'mDQ�[�����T��x �e�S6��Ձ�Zw�s
g��,��v���ek�d���dI&{xK�d�h9�w�z���i���7Y�X�>��K���Ml�h�k��@�-�V��b3#s��q�K�LC��G�g�{<1�ND*3�h\A��L���\��/��"�e�pjjր_%�j8�B�S]_��s��ȏ$R����Xi��@Y���9LQ�������KNT�)�|��ز�?z�잰��������G8����2$;��{C��U�˓ȋ�@�����MG�n�V�~9�̩&y�[p�/8���_oC+�\�N��/s7(t�'9��mc�}�t�S<��cnv��-1���_U����i�q�S&�^�SHӏ�-F����%;��G���6�+��\�aX�����31ӏ�������%��F�a#,�4��/"߉!�*��.�HQձiQyϜ�J&`Fm�AO�KxJ���ۓN�W�	mҚ�� ��m�M/G�5q�h�18�ʤ����,��cXÅ7�9�߃���n�v�d�v�D{�����"�3V�Ř�5j��x�T����U:�8���gm�2�� �����\+���4�.W~ �z�\5z��0i�RB٩�lL���f��$�_H�E�H{<�9=@��먠)U:f�����Ш��@�u�U~��2]�����;�8Š����7�xG�PU�Z��&��V�)�o$���{�C��mph�1Ȗ.�w5�#�D���mF�u�������O���l�0�دZB��K��ʎE	�/�«�O��U'u�Ʒ���4P��[�z�_qSC�9�"�AtJ;��G)��d�_ZaNeЮ>g��}'��`-�Ś8h9r;1޵�}���-��4���Isp*�z�x�J���D�ޮ�K�6����U�عlJ�}6it��� �Ob.74(�
תR�Am^B�b��^��QO"9D]<g��}F~nj	K���˟�ڼ׾Dy��Ev�s�df:��=�#o��տ`�5����˚����b����\x&"z���x^O�~��8+�s�V���=�\��?N'_��A/p�ڔ.SK�5�.�Fx$�j9*�фB��S*b�7{��5���SP|��o�.��6�I]�& l+�5_)zmj��Q�@(�� �&��D�Vn*�Fb��j�eƘa�l��=�lx�c.�S0��
���j[/��˶y���1$d�O,4os��k<�
�1;�]Cj۸`�� ��o�h����p͐����"P���[/��l �Ģ`8\��R�9���р�U�?����1����;��}�<�i��[qph��j�"W0�uG�u�Ǿb�v8B{�{Ͻ�B�[U(Q�+���X��>%kx���\>b2`�d�2���z�w
L��旫Ѣ*�Y�N�M�xi:�1��Q�3��}n�<�|�E2���T��·[K�g�t�&��
�J���������фy7���P��s��ˊ�5��������!�e�!(�e|�'`A���m����֪q�n�t&j�D&f^�eLT(yM�����迬7.�	�oo ����-��<�w���K �Wv���X��Z��X�Ng���@HJ�;X�y��������t��|\��F��N���R�9WN~]>rwS���6������\V��\��I\��� �b�'�����81��6�ٺ��YQ�CqM�����߅��r���}	����s&!�Dd�c6��Ύ��ب��r\���Z0�fL����� � �z����^��� I�D�	?�J�IĮcD��a�B%��zu��T�y��a���v�P��t6��.I�����k�$�ռ8��1�غ$���c�o�{T;�-�2f��r�Y��}�0I��{{�X��b��n�N}EE�ߦÖKP7p����<]��f����0�C��EjGp��Oj��� ��+�!��ġ��B�����jџ�>�QA"55���T�fL�*1^Sl�2בʙ�5�&�����8�|w����f4����dռV�i&,����hr&�/�	�?%��|��n6#f��1��T��-�ߢ���S J�����ҟ�k�n;�� r�iZLd�x���uj��L��k��C8/M�}�I)��e*�&��G����jV:�65�	
u��l�q�CS�
(�d��p.���d]����v��y���[�X:�J�lw�͊�X%!��ĜVd�����'���7k����ɓ��N�UP���k�}�t����Ґ�W.Ձ� ^g�	�k~�p��=!�mwY8�&���T��n�c�R�:�Q���Z��XاMU�67����QՓS�J��i�Fv�oЈ
���y�6�`l;�7��yEl��I>��b��2h�Iv��_ l����g'���g���L0�n�W{I�_�0=o	�ųONt��6{����V�6g��$x�����Q�bc�2�L���h��2g�2�!�
�%X������U��!�I `�F2XY��8�H��#ᣣ��_w`&���pdk���4"���X��OU�%��w*⫰J�?I��k���T5O�l��D�y'T�7�/�ȓ��#2|X�7`A&n�� ��U�0�Vw�K�n��u���#��h��[H١�r���Y�>�bYH.��x;sk//Gt��,�(��u�"�,���j�9��Cd�W�	P���m�~�S )=T�����0�Z�+�?����O��pn%������pm��v|�~j=��[�4̌_��u�����ƍ��*����$��nO�p��'a?΀����B���G���e��G�Z9łk"]8*d ?�ĕ����J	]�C~�\������X�J%ǳr�x��KϟJ��딃dpr�.�*ըY�f].�~I�9ͤ�eKJ�*�ɑ���/�E9�����A�s.D���jÅq�&��T�/ŵ�	"��Q�������h��|�a��wd�m�	7���ss�>��DK�8e!�G�����<K��(+'8QgFXw�*��j�ߑk���D-��G����3:K������t�b>SEXP2�_�iB�@:a�0o�[6��ڞ&^y�i3�oj�j}������?�|&]� ��
�8/1�^p��-
�/���Tw��	4K�0����H
� ~���k5�������D������)���~��"93x�Y:��Z͍/}�{�U��bX��ֆ�C&t�n���E�¸�~��7��(Z#(m��g,7>��C������x+Z�f���1M�-9(?�os2�sG����~��-���x}�3��B3X��*����;F<Tn^ЛK�33���tK#�%���<��������a����/�!��_�pS�d���^���)<ץ���c���-�Z6`ҶFg�BqW��]�Y��o�P*��e�u>އ�A7�3�����?v_���ut^0`yjt���)_�L�5~ٺO�7�~`�t���r�M?91�X�H[YVC9	&��Ke[�'Ay@v�:�5�4��}#p����ia�1�a�f�Y<���lV[ɸ>�������2���d�X������.c��p��
�Sl�����tOK7���u�'�;`(߭H�<�k����~�����Ͳ��+���k0��q�*�l���P��3���7`�GFI�k���_VN��PЊ�z�;��v��� ���r!I��z�{5��}��-��GJ����y�6��!��V�͢�MC�m�^�A]K"�1A]
�s�@�va�_])?���%;�&��� "ݖ�~�C#��]�*Ĝ�e)�=]dԀ�2Ć+<z��g��,kb-�,+LI�f��]�Z��C��X��r6�548ckgBg.F�~����z۶E �w3{�{�[.�J�
k������"}�\J-&Y\nӡ� ˹3F�b�9!��>}��CJ}XlxV64EB    fa00    2aa0N����[k��!�H^ ��U�R��=k�
�X@c��v��~x*�B��-�V%
m�0d�Kj����qNj�����hK��J"������D��Y��El�T���7�������z}7VK�"��H��m���l�I�u���10�ĆIGָE��҇L�J�C�Q[ j/,�cZ-"ü�IM�.���ПRO��yЊ�Mx�7R�Y���ͥ��븥���X�0{�zFt�J�m���&��>�r ��^�!3�VGCơ�����s����E�ge�����JZ��C����T���'�5U/��ן@O��.j��߷a����G	4������%<j�c�9q&�9h���N�|̊r-x�;�s�Ͱ��Q�
E�L�k#-�{�Qqw�V��|5��dQ���&�Vm�����9#Ky�Pi���ˋ1@�B.`��Z7Sj� PQ|?2�F�3��i���z�r��:�no��H$���M�?�Q����d�䭇莐	����M1��B	Iz�P�����O���&gM#�%�<�Xݰ��hf�2��Bk2�Y�J�!>�,�V���v���E��ۑ��T�S��9(�
�N�I${PE�x�浢
�dh)m2�$=�[�:���z֮ս7�9�Ơh�G=,Ñ!I.W�Y�.Ri���e�BA����Gx�<���!���7�����Z���u����܃&Xg�#OK���Zl7��R�D�y��k�%�s&M�����`#U���a9O�P�d�3�/?�"@>Gd���V�ֶ]%���F�Wox���,��c+o�#D�Zv3�â��\.����P�R�t&�P=����(���%{�
`H��P����GA54Z-��3�63)����<!�1���Y?xj��n��O��\׮�8H�y�3�%aG���V��_���RL{�?�Vy��;�P�,6����i�u�FBš���
�E�@=�9K�r���2�̠���?p5Z�:��P��܋�:���ed���Ƈ�# ̖������r��R�@�a����4c���-�)d�赵h�ј�1��9�̢��E�7]0�k]��.��ÁR�
�be�D��ҟuq$���Y3�X^�9�r��+-TҍC�3AHP���,�a^O�y�� ��4�۟�z�B�Fk�V�j%!T<3R�q�����S0X��	>�W�z�c�RS����)���g�c�����mh)L~�r�[�f���+�{�����-e��gL��˖2~��iXbR���I��C5h��9���:m�% �N�� *��-Z� @D�p�]�z�V���4M6��%��'� ��ި� f�I�u�8�W�ܕ0��V�X�}v��|@�j$0����f��8D`���k�c4�|l
7r:��p(����úN�ѕ�F�8cϰ�dW�طi������`���P�a������J%ݰ2�
�����Y-BT���a�p������7��8��;�j��ҝŷ�il./�"��@?��9�e&�!����8XC}�a����=����
�}����J79I�H&C�%Ų�u��V�`}e-.C# .��]ef*�8ύpA��`�L�8	R�_���^�x:g�P�a��HK;�ᄂ������4g�]g��x�2��&j>5*��*O��r�0���ʝ���� ��`~��X��j����͜����9�����	��YO�ծ}K�� �o�ß���K�[]&W0��zM�q��%�i��Va�� fL0ݎm�D���>8Ţ~�����jTy��� ���Kc��E�m�՟�?6k����}��A��4�����=*Լ���͡oPB@ac;��@�� ��Z*ul�oeT,|S��sY`�@�h8��(�J�W���Z�2�<�y~�f�Ml�ō��V���}��Zep:�T�(��nO�f��\�r�^����d�1�4����>!�B-�FYd=P���D�k�̓95�"L��ӝ=���~�r.68�)q?��,_�@��`'�ӕ�nb��U����$�!h���U3�>mw�k�tP_IK���.o�en�G�@]!��1��`�M�� � n~?���0+/�ǱV���L,k�``{�.������M�PN<���4���>H��t/#Q����Qc�u���M��O�']��o�K���!�(y&I'��z�ҖPd	����!�%���.�0X�Z��)V�ho�B�6�*�������ꀘ!F�#B���tڑg���v�JZϺ7~����������m�^�~��;Da��/��:pX)f�~�[n�O��⣳��I�՝��6<k}9�W0�)�B<]{FN��,����}�1��ǂ�����̗��:K� Lw�?�ߔ-J.�S1�E%P���~ܺ60?B=DB������R�WTr�>��K�?#�ciJ�V&JH�v�xg��_�{-��n�a�L�Ug)�s#�Z[O�<�at+r������"nZ?>T�U��L_��_^e��4͵��O�����.e�AWp�׉�|�IZ�}�}�DF�H7
w��kq���IGag% ��u�4��?�x���7 �����Ugq�m��t��!���O�Bz*�Y�������Һ�����������N�=r8��49�n� J�#�ߨ�fQ��9Y�t�'�zm�<~Z��3}-��W�+d��y47B��Acj[P�	1�t�u6)0��P07�(��u�3~a/n+W!چ� �ڜ�`�_o6UR�U`���\=�POv�Y 3V��UCwH�̞�	�n2���t�1_�È���yܾ�	ƞ'L#2��qO֋���.��Y�B�]'"v�&|E�"k¸���4�0J����!���w�
dq5VK,]h��᭛C/=w!0|�c���cr@B�Mr_�!�Y���9��0-�^.��O����ci!�۟_�<A����M�ߡ%Fc���3!,>�&-j�[�+���=�]��p�/�'����➞��i���`�y���FK'�m*.$��3{s��C�4��#�OQ��|�/��ƽ`��,�W6��t�Z�o�L��,����U��킸j;��+J��7��a���`<��۽uC3��<>���΅)P�x�ꌄHf�Z���-HPtԏy�X_�iW�?�<珈ĩx^��v�u&m�	�D	����p	ji�� �8��Ļ'����	�vC��?�J,�1�\c�1$����Y�|7���$ܷ��Q��
��D�/I
��F0�9�q�C��YO����bi��M�{R�W ��T���e_@(�uçr-�~�Nj���c��i���Q<i�b+>�2i��x���hugj�ˇ��-�\����'5�CQRp��
%B�xC�[!�۰?�|�D3�0�l�K��YLpHV���&,`�;�rxQ��5��r�Ҿ�N5����Z\O@՛Έ�Y=�͙$,��[Ha��Eڐ cb���1��џr�j����&�w�{틫�H�`�ʍ������8UG��,O$Y[��*1[`-��*������
�	� ���z���enlD:�;��,;xG�;Yh��8+���.P��X���:����+5��3������q5���7|��QM���X�w��XwȠЎ����H����XХ���Yl�R�
�M|X*F���ו-��L<����m\9�XPM�^6�S����-��P̺�$&1���XH?���ͯO���w9*�i���x�@�w�8_(�aD6��������'���Ej�\	OX�i���Zb�F�ѻ&��/m�e�T[=������U�'H�B}����'�����-1��إ���3T��{����V�
����M�V�R�� �\�b)�����S?����O��|����c�I�@DŒg��Bv*0�8j�q�)��/ݧ�F�䥉d]d���(7@�=V���\��y�o�h�l�y�Ҽ��{��&�-^bw��Gp����%$c����љ�y�t���pB�Ivn�-��uO�F;�I���x��\�q�|ޢ��O���%l��n�P����!�1�!�TNKd #�!�%c��H�������o��W�14�MNLf�$4Xn�O�7'
4���]��)�S��5���D*͛Ź�Xm������4�)�r��i9sH��zV���M���ey����d��~|�1sЙ��a�ɪ�#-��3�ݭ7!Q��Kp���{����vt�t����г�s�L���d`���ȓύ�d���"� j!۞�%�/1���ˋX����0�Np�����ZB��m��mM+�@D����G��P1���)��-�ǯ�ث�-��}���,��w�>۝����)��������O��¦�|����"Z�8���/��e�J�@T7�-�S���噀��|���s.�C�����H����7��Tk1����G��o�^�����b��:/����F�cLC��+�{(I�\�[�H�å�v���.S��N��V����W��;5�u�xe^��
M�ZoV'H�!��O2�Q&���ݰ����B�=��
�	�$,(z9	Ws���~�1Ӝ�2<�E�.�n׌��K*����::��R�Đ�tJ��̯�*YqxYW� z�ȦI.)*�t��ә]6�/���H�����l����y��2	��r�}�a�d����;w��Nj-��r@�4���ڠS�ȿ�D�k�C
�N��Z���Lʴ�T�ғ.6T���9��u�l��[d��̑��3�����g���~���o9y�\d�l�"G~���N�-+��6&NA�3�I�m�z���`�(h2y�$z��"\�cs\�vJ�D�T�/��H��+|W��_�f�Hl��'3�&|E�w�l~g�t2q���iA���b�8\����[	N��Ap��1���t��lf�>�L�4x����.xD��6�^��?�i�s��4c�fw}����Yq�{ˍ��s<�~�����{~�j�-�W��M4�X+ �e/�v��)K��M�b����8�Z�8�:��\+��!�˜�r�B��P��R����ʹz��6��q�3C�����|%̉��H=���o�f^J^��RQ�X`�^�D' + #����^j	��2bFUS��M��
0��۷(��i;��5��h�ٟ8ha֯0g}z����n�#���<w��^]b���rh����hR�uel��Jz͹_('&2�d�.Gea��oÝ���5��7.<�YVq�y˳ӌ��j<��D�GP8�����6�΂���6����-����Z/��Q��jxB3Dc���:��w��=Ҋ�h��%����)�j�֏���KBߕ>EU~]�!��3�S^�m��j?
�ܟ��eR	�����l���6�2Ee*g]�s�w;�󐫆��jQ4zf��S�D�JrW�dN�*v���"OH�R���6����7XD.K�����]��2�
P	Ťs�ͺ�7�;#�d|_�}h�G;�[kT�U(U��&7�%�� ��1��~1�h*�?�B7(��.X��m
���'�n�왷�
�l+Y�
2u��1����c�.R�_H������`<�	p0O�EE��:�0Ϳ�o��fXg���zAgΉ��2q��{���;н��կ�~I�-�I�8��/��C�A��m\�]1<3��AO}��M�*� ��S���s#�_qjӶԖ��'_��`N �m�J����Y�,%��t/:���3�ڊW��qF<6��3!9��jVNꛡôW����I`�_9�_�{�ctK:o
��ܜO�,�*u3(�Y���q*���+�[�^�Qd>ʎM1e5�� Б��WN{ihe��~Ҏg����m���|Fh2(���z�4b[I4�����d,*���:��e�U�cġW�89GO �^Y#^���& �x �˰?������EG�r�-T:����0T���x~��n2�k���'�>�IS�����)PEK�ڧ�b�*�<�%��f���N��*��._�g4<��tc�)�n�q��0�1Z�Z��î[;#r�k5+	���"�\� �yFk�,A�Ğ�t�)�am�3G�e�w�y��e��"�epAp��C�嚂l�ӆm�v����	��^�b�^c�u#�9@2p�kw�o!y�B�Ѷ
-Y�]���%��]��fhH�E�v�g��shA<�ځ�5Ɋ����4�E�0�9v��'��OQ�oV_+���.'�}pO,���B�m�u
�c�)j����=U_��]��x���@�|��|�V
�8o�̨���I`ҔUlP��۠W�ΗA	�� � �_8�7S~'>�����&c� �E�Ԯ�����NG��o���[�vXdz^|��
�^�����C����d����{ ȜлO�����}����U@����^ԫ��Mu�ێ���yp���1��v�ze�x=P��&�8���BV���v4����@z2��o�����i��H����^ߩa�{��i}�Œ���>�j�i|ڃ�j-00�/C�א�{�1@n�a���bYm9��-����W�I�t4=��Q�=���#~��,��#�r���-n2��6��U(�bY������ť�7�QZe���cy���.1'�lЩ�?�k ���`�wX�qi��*%��=��
��I�,6����_�V�/7;,�7�_�h�:����ꛎ|0]c�n��w�I�%�EV��Y%䮍�h��^r2���2+��-ʒ����d{��_�n�N�UkFt���BM }��Y|���9x�-�؂�_C�/e��8&ݏ��N�4.E���v
۴�=ճ!��G視�+req�O��@�u���*6g��%�E�"5@ a�"��b���<���qJ�Wĭ��(v�U����h��+΁w��<(:��k��|Ý��	SK �%�|���y�? ��e�˛�K(�CQ�q!8.�W��+�߻�s
y>%/��ݤz���l�b���O��������%�n!;������3���,�ض]��@q���`z0v���S�rG�]��k9\fdb�:R:e.s+�����WK�x7Im�c�|����O�9-Z�B3��f,����*�9��cj��cي�/��������K����[51�����*����;'|nu�:k���0�.�$�2���+T�I :�˞���ͮ�W=z0��H��(+��o(y�\��4��W�[#��?���:L(�w��x��] �ۉ�N��/<�%mΐ;Վ�~��C�<����jL)����F�8�s[	�[}]Qso����E��5�87�+q�J:B��((]��� 6|�����|��)����L8F䵩lp~���rr�%ٵiE��%�ze��)h���p=s�4v��o�i?Ȱ���&��r�R'ד>8����)��&����M<�A���G�X"F��J.)�ە�+��]S:��Mz�Mr/�������rHf�8�ݱ$�ݺ|�i���7K�;J3�`��'����z�;u5sk�Iy�x�B��t�BUZ�����4�`0
�ͺ?d�����g"|�D��yk���,��CW�U�$��W�mkd�o�R)��3��g��o*p/�F%rL���W���x�-X����1��F���[��e��o���6�OǬ �'��@��ya"�@0�+>��StP�����p�A|l���uA�^�n��6���F]5)�4��T�i֠�=��3�T?v�C�7���[s��t�����""*��q��q������2��72�")*�D k�����9���qs�u;�<�P8�oOK�^M�	Ԛ�N�V��x���[y`޵�g�D2?a��G���b����sUU�6���ufx��9���e�'��R�o0-u��kķ���4�D� ��
/����x�Y{��Y��S��{���8H�
-+�*��JӜ�j��\��w$E�de�4�sI覜�1�V���v���_�[hvD `��-�})/�WY�L��I�G�DJ��v4��Q+�#��J%%�h↰��P�%��/�+&F��݋�R�āL\Y� 2��xFo9�x��@5������~��7��1h{�7��T&P��nգ~:�h�<$O��,�N�F$T������Y�G�X��r��79U�Q�0O�v՗�ڴS�zY�x�����I�xN�|F�Æ�[��AQ����Tk�=(��-�5�X��}F�ks��G �(eDV��?+.]�aB��5��;�~��NP�#_%����#�7��k]g�I|�s'~��bޑW��Oݧ�!�&%��e=?��O�\�b�颜��0k�Q,b����}�w����fop�����d\��'sx-��|Kt�=gYt�0,/5��؜���:�fKcPƤ�o��� �e�ig�����i��2�nJ��G��(�5g��o���Ӏ��wt�~1����.��f���-:�i�
Hn\]t-���e3˲@jv��,{���Xs���,�d�2<H-v�|����e�uh��+m`D�wȻ����R�=���b�a�Ӕ�6�3�^i �b2&n>��X[���4��l?�a��-�ab�>۳��~�D|Pok;N�5��`]��|t�0U�ٮ�B�rX}*�6�\��!v�xY�5��Jx���(��Q
�tK֎�@�<2��Zg�A��Ns��t�ezEz�Zh'�����SF7�S��]�I4{�*�Gu]9У���A�^Z�����c�ޙ�+
`ʪ}�q(�-9�m����h�Eۈ��L�kR5�ۃy'5��<��Zr�Ξ���~�xFg�Aqm�}�<k��|24��i����B�4���3k+�����\�n.�Yi�ɪj\�.oX+,JÓﭻ�u;P[�$Aޖ �l��@� �|�9���!GZ�Ҥ�]X���FR�@���:��O���a}@>����|�!�s
� O�q��CC��v�M����̱����ǝ]J`?IⳂg��[0i��=�[�O��#Hb���Z"��3 �t��m��1S�j<+��0��D�G��Ӆ`�m�'#�Lj�`��OP*Z�Ʀ*0�݇4ށ��3�����4�7��Ԓ���9��a`n" z�+3�Lz�i�l�Kvj�]yv
�b�E_�Ezw5[����%���Ux��ݏ3��5܂9��!M8 K4��Cg�l�z�0�##M��������_L%�Z���Ȍ�3�l���R�t}Zc}8���}�=�}�Eb�����~�ſX`�wd} gd��)w�Wق�f/A�]+<��L1rl,L멾B�dV<�DvH��*��?Ý�q>|���k��h4�Ci�|ʅ�:"�I��;m:yһ׵�/9:9��D���l
��,^^�`?V A�Up�A�m5<[��llA�?��іһ�(K*^���1Oe�X3V�a˝�Sx�u}tW�O���`��RA�^�l��q��c�h��e{Ox
�cd�ûv���a��.`�HsZ�Ӝ �t�삒:b���Ŋ������e�& 3��5C�K��OVx�ir ���ׅ�[��S����D�x���e����:��z,�ѝ���ĎKm\eg�|����訿.no'��}����F"��B�r`�t��#O/�i�b�6T���n��}y�>�����+��q��uN$��ϧ~+XH����®|�8���H6�cX��߽'��Q� �ƽ�7����U�1$��q.���+�kG}�~�)^+��G�΢3/�
o
�dr_��ެ��ЫCS���t���L��\t�w�SST˹W����1EQ&�\� ��LF�6X�=]��$r�3���)�;LM�X�
�Y��:m� ��dԳ#�k+͔h�����U� �'1O=������g-���VB9���ګS��i�/:.\�6�,��p4u���6��%���x�Ѩ[��o���z�r��*Z �&\e�%��f�v=ص�n7�"�]���=�w��"�3����������	��r��K`�Z1�Yx�P�m�|V'������&&��$����>,��	�2P�䅳�4�A���W�k�E1�z���h-���>ӡ���[�1�o���rs\o��A5�_���{�X�[��դ�S'2���L���>��Ѡ�� (�
c�,����h]�����c���Y`z�D3�:&߆�|��3{0�љ=?�}m���0bO�[Bl��|��`�k&���t�:-���Bzw,�Ԣ�D���	�]2��Ϯ ��n3�}��ק_�iM$^�l�J;S�Q	CÄ�ک��X+0�16:	�5�$|�A|���R����B��=b:(#�1.�2%X��l� wh�J�W�4���𣪞�[��=�lь!=�u3�ޔ�ne\oO�e� ��RdA+O�8ۤ`�!w �؊�����ݴqu�p��n�_�b�~�Jw����[��q�%G@+,��yK
��#rx�Ϣ�PI�|�ļn�>�:^0�)F*�Gh�y?��9�y�U�E
,��x��f��[8��:P�j��R��S'&��PD��7��bB�<�q.='�x�����MٶX-���UX��
u��������� �fk�'@�-��a�=�yyސ�����d0L(?�-��:n=K}��Vv�f�y��Wx�\�80��C�xgC�k{@�RcF�K��^�Z�(�o�jx���r�u{̳]�U\$?�L��\��	e�N�:sˮ?XlxV64EB    fa00    2750��5K�r:p�J�:�0�0�-	vFʑ�
��l�HD�x�g�l�_p�u�>.�����sh�~"�����	sV���5� �t�|`��'0�1a�y\�#x����� 0mޜ\eG�УV���P���ި���MWh�S�1����eW#��R��7<E����9x5�)��a�u�&�[��u��#��p*�lr�(I�Qbg���]�)ZQ��d�<	�/�N3-\��ă+U���]�8���Bz�fP�H:�/k.�w;ak��p���5P��p;4�Ejo4�s)����(D�=Z�p�sK_Wy<W`Nq�0�pɛ�	S�`X��>�\�L�c�����w7*<�d��!�od�����m�g|X/\�~gM��2ѩ�ʎjS������6�j�@+�c"�k�N�[0y�.;�Wmm>wm�^ز��G�}�	������q�A �"cÇ���*VK퇸]`�. �,]����Vr��sj�׋C.�D1N`r���8�*����Uǔ�s_�x�"":�!<h[��������:^o|�*�t�yN��d�|�2�4/�] [�3v�Ԡ��Dw�$�1�2��e[�����w�R׮�E ���O39�
������>߯Nҫ����ʓ����%0�s��P��|F�4`^p��>��s�Wf/�\����_j%�`-���xj-�c�׽#�=;jH"I����g����9'dy&0x�H�E������X��!�2��F#	P�\qfC�н�H)i �*�A����N)"�\���s��!�x.J�ן�N33���#|���j�9�)��f]nԿ������c[���	�Zٱ��C�7���¹?�^C�	Dera�m��0j�Ag���2f��t��NψChVpұ�p�o#�@t�~���1M]%n�7T:���l��6����N)iZ5�-d�K�9����>����"����c-7=�&Y�$DN:��X��caR��|7F�B�l,�y�_z)�rq���G�j�|)X3� h��YHe�XJx+-������+k��"�݅�����9pq�nl:�k�qNPԘc��@��<]��-����,`j �<G�L��l��#Md�*{W���WJ Łg6�x�۪NL%3҂�.�4a9���[����\a�<�`�S*�� ����$+a�M���Ja�0�O �#V/O��UX�v�?��9O�I��V��ʳ��L�^~����*���!T��9^ΓP�Eh�p�K�],Y���jHp	�X�8��#��q�Zk��a���3�T�x�>jS��p)χƋ�&3A���U�^��R�p ��[��ɡ��P����9��>}��Q�����V���;3Լ���)'j@Z���}�5��m{�V�X��a<�,8��Ǹ�{h�i���[���0̰�E�r�`NdA.�_����`���>��p�J�t��[�=���ƃ䜖tS�䝫���)}����W����0L�_F+Y�w�'e0_�$m���|;�R�<�aó���E��عUh�PAʢ�0���#]A$Mdl�2�c�Z�`�l���T,X�
]!GE`N	�O_{�������\�(��aB\�jq$�q�����Hy`X�0r�y[�1I��i`�7L?_pD�hom	>--���,��	��jr˗�j?��fRT�*;�qx��zve����Et�uJC~��$��qwx�d�DWD�آ���b��T:��v��x�N8N�d^��y���N��lI��&a�%�\Ӝ�9���C]��9*]^gBE����z�1M�tIgz`��TYb�k�O.�c�i����P��[)� �%(>��Ѽ�6vKf=�FV�|���f�J��{hp��]�FϜ:���\IZ��t�\��XT��pX����#�^��������n!	\�9j��|h�{n"1r�e�6�ؓ><��2(���g���҅�����6�?�-� (����u���Z(���u!��cI�ú���
V���ju���NDBp�*ZP�Ŧ��(o���&�새�B�h�'�K(�b�`%�3[���{�cqS5�и6�|��F����)vfO�_X�.pu�N�';��>Nq��;$K��_�7�@��~;���}a܂�E�7Gmp�Y��&���/�W,2��������)g���MNy���8�p<ͷE�}w�%$��x�%?
���.�F�CTܳ���"�P���R,����8��� �1��,|�����֌�8	f���tCW{�&]�!l�8h/2Ar{i2���).xá�&�:����3٤�����l�=s0�:,���3�R��Q��W��RbG�N�9���8A�J:	L�@n�{�v��=���=,g��0bU�7l��A�)�/�j[c9�����G���.��~p�%I��)�#�J���ە`2��R�V��w���K�G�����Ѣ��3%��h]������t�XiVY�Y������m�ed
醧�(;�M<�g^|㉖[��ȴ���,/�Y����BJ�ɟt+���%��I�3H���l�עa��k�-
��;}B%��i�IMܒ�_�rm
��Cfq�'h+S��Kݔ�.��H��sO�C��I�/9�%�y�:JFC̳�~��Z�[���c������.�HE��([Rxe��^�(�?1vjH3$ǃ,�r	A���(E�U#���D ��t?�!� ���8ɂ+.E>
F_K��N�e�"��/�HFUy�a�SQQ�x�O��[�l�C��}�o��t�˪�Pl)#>���s���7^B���^���o ؕb���B���z~�>MW�A�I06�k�09+�~��X�Ʌ�5�[��IA�QgJ`���.4j�ʜn�Â��:��&�u$S݇�kG6���m�夠V��ϗ�v���8%!)W�?&�;!0��yGZ�(<(�V��{-�}�v�U*��dѺ�����g'W&8��%�ЋKT-
��#%}[c�a�ǠgYii���v#��*���G��iYn߼���i���7���)=<#ꬅ�+@v*W�9�]��m֋"R�cva�䕬�O~��6UeD?<�1��>N��zϼ�ˀS/�s5'�����S�{qq�����-���-��M�	Xt���I�M)����|��ş��`>������F3�~�eZ?����gY��"&���ՂWP�����,�+��Q�X��鼧i�b\K�̲O�g�@}:BP_}���n�xpX�}3�T�9�i��E+��^T���9ѥ�8a�|������=Q�՚q�$�ćׁ'C@��&Zdd,b�.�O>�I�b�[���d���܀ E �����W�J	|��9䡳�.�vpS �h��*kF���4\e	s�H�`��FU���#!/�@X�!�s
'J5��O�M<��|�jU����d��v��I����DG��0�=Y ���1پ��2: �R�*R�0��Z���U��}�9�k�Y�Rxb^tf��Y6���Y��F�(G⒡���<����:�k�3<��@$n9�s�JB�mZd�]yЅyx�7n!a�Uˡh��n��j2t�ţ�_G�V���DA�)'��u6����ޖ���FQ3Ky�_�6��l�$ĉs򑆟��}������)=��ƙ��^�luˬ�ц@#�Q�wWv��#�Ms�9�'��5�w��g�x��c�ˏ�I>�о�M-x��j�䯋ep�	�V�n����*��۞���B��m�B��G �-��]=M��̦�-���^���IđD��Į�[���Hc�qO��d�n��*�N��B�%�/���$�2�s�
�E�������|����d���ZOR�2��`ِ ��G��ȶ��]Ӈ"�Ir)��;�/�����ʮkX5�47�z9�ٌ��3���WomO��= �׼���7w��V2�8�Ȝ�e����@nu4y3�ug#}��=�@c���̉�&��띏�|4�o�d�1���7�n��e\\��$�6Q�0q�~n�l]y���@������y�1�fnu���V�	'����wi�\�6n7��w�AZ�.پ��!+K�C�w�P�&�$pm8�W����N��L��26������Q(��0�����)��[�o�@y�P�i�)r�}��h˾-�e�I4S>(��qԮ��jܭ�t[�N�@.a(����];������PQ� ��}��S�;ُ�m���h�Ş��`UGI��&\��=�y���-l���-}y�{G���"��ɫl���I1�{�b�1��/��s@ç�9�*�0����s�Z,���v�>�m�I�
i�7�=�����_sMh2<��e�À)�Vp�'m����X����3�e�܁}���Kx�Ӷ{I:j\�(#����^[��2�d8
�nu���݅~������;��O���M���8�mϭT3����pV�*5zl�?��h�Ю�l$4
;��)�Җ���<��|m|J�X�4�2�ƉK{a �˚2���5pf�]�%�浈�L��U��$��+����25��8�4�W��L1�:h���Y�Ѕʘ�b�t��HƓ_�����/�3>�b+ONe�"pNu]�����ȡ!��@�rcC'�KA�1�)�_�8�	I�<�Q}5s�������V+�G���ި�Sb�YU�e���E*y���B8�|/�[i��ؙFb����S������P$r�^ۅ��]&������!��t�B\�S(Idꗭ�P� ,jƃS��d��!*|S���� iz�}����<il��[P���ǔ��X��>�|eЈ�lx��ik"��(�M+�B�kt���BQe�}�U�g��=���?�LX*��ާ�w=wE�>��I5e�7�㎑F�~�T�xkAm�ZŌ���1�QЧ�[xXH���."g��b�%M�qo|���LE������/��`��b}��A�"�H�n7:�"�,	<�p4��V�C}Q��X���8%�t/R{�`S�m~Y>�H���
u��_�O�ɂ&���Č${K*%������o��p��kh8���-��k�X=�'���|H5� �"���N|T�ʧI�]q;i:�nG�R��h�L�VXܲ5��ߜ=Gt�!���ZS�?��sΗdJ3�0���0l�>>|+WR�� �	����
�B�v+$��"�%<[�%t!�q�#ٴ��v5���g�J�8�ʩ���,��P�a��)���ϟWl@�_��#���4
Vx9߳��a�sl��b|�����b3�3{����l�-e�<RgRKi�.f�L�R5n$�I�*���	MG<�!�̾�dj�;�zu���ᕞ���u��Od_?�z
XW��4c�C� &�6����T@"�5��#.�D��?���[�:�Z�7��\�!&��D�e�{��R趒�JL
�L��"�0��0[Ӕ�V)B�2���9w����y?��3盻E�;�k �|p���宖�M�+4�Y�L:��3eYK���ϱ�2����(���$Cȃ+�v�h�ѺJ�r�C2D����LHm >�r t�r�S����T%'��A_�N˹J@H���Oj��I�~'D|�mk�MU	�$9D��IMA��#c���M��H�川����e둜3_H](��i��4H`V0q���ŭt�/�Gz-،����\1�@/�L��Ռ�:�_�e��Lμ�r��?n��5&��k�v@1v��J����Yë~��zt�G�g�����X�]Z�aCG>��7vZ�b/s|�&��@�v�$��f_Gc���.!5W��bL�#�uTk����@)!�@��e"�j�7�̫`�U�A[��y@�o��l׶)���)��s���������ز!���,��M)���I�%����ؽt�ta�3Хu�O8�9<Q@8T)0�k���i��M[���Tk�B���}kA����ЙX"��H�lr+�as���."�S�+��^=1��W#3��M�� ����;��d�'Y2q�'�z�,?�݆#��G��Za�i�O��͒)���/K�/,B�~���^]�ɽ�IU5������� ��&�{&����O?�!X�N���j
��t<��O��ҧt�,s����bt���Щ1��2�Fw�<T��A?�����J=p���kWU	�׀�4�X!��9�����oG�2��
�L�;̈́�8�A!�+M�Pg��qd@��*vܰ��`����4,Ey�*}�Z�� �3��ή��Q6�&�?��M�A�
8��z����:���W���MמM�|�Q������~�q��_V��/u\~������s�id����k#�q/�]�@�<�����|�y�9g(kک�eiF�袹?M��H����O�S�s�\���8����Qs��P$�M�tN�2��ʽ��N�*�=j��mF�$�'�����T�4gz�0������P�8��M :�J��RSZ���h����w��L� ���ga��1}�h����\;,C@�7�ՑapFrD(=b+PXF�W�c {��	<ip�����1��I�+�k�ai�z\�Y���E�s��͈�Sz���,���%]���1�d�����h�C��"m�"_���B뤹kLi�t�j��v�����FʇZ���]���I����._��R�)�_��r��a��3d��v����a�ɘ��+Aߚ���DK���0�~��Е"۽{D���0��;�6��
��Z1�~��W|��h��:]�ۻi�US4���h�}J�8��>�+k�*�-㊼>ܵm���Ҁ�v�^�E߂%� -Ӧ�_�Phc-tC٫r�ܑ֙D����F��!ѫ���TaP8��J/�5�$����RgE�����"@r6Zw)|�F1yJ��oo��ݓ�0����Hx����FiB��K��D�?ڵ�4@���H�y�N�59;_[u�W9p*��#��MM<�r*��Ԣ�L�ߓ|+�8��ݠH�|�lA�ȶ��(#�W���y[@��"E4$_:K�~����'�<9g�.�l�u���̿-��w�39]��v{���(ey$
�1�CK��87�7�d�q�X3�����Eh�H*�{ ��'��V�{̕f�<��^�/���n��M�iT4�3�����s��g4��C� �O�RF����w`D,��܆xI�;��.�C?�N�,M�7�ͳ�1���S�7�Tٞѱ����F5���#v-�
#�B=v�E�r/�:�X��t�7>AE����t7��{��s��ھwU3VH��5����˩���F���-�"�".��̖�C̪s�*!;��Ӿ|=�50��Q�Wf�m����%SV�Jh�b��b6!}yuA$�V�G�7m����g�T������Wd��$�t�>�ᑛ;����٥z�g@���5�J��՝�W��\�R,�w���7v��ĸ�,�W�/�`��e���'I%<�1�#En_��Sa�^5��<�aB5W�Aj�![�;�\plW�_�k��+���� 6h4�4��q1q��nFG�_>BA���ΘUK2ǧK|�w��0sk�8�]�Sl�E!��!:&m>�ю|QP�U�H!�i���ıC�v)(�*���̕j쳻�\��o�� Ww�*@F���V�S��rk���L��=[d��	ϝ4<)(�K� ��zb�S��R֪�\V̵�������ħ����x^�8��˾�`�3�vB�:E^�:x���%f(����4�s��-�8�;�Ӿ�ʱl�(+hZOa����Nl����v�l}��jjI]t /8��H��:rº ح���V��)����;f����?��YA�o.�I�r�U� `rL�n����m0�����P���B�GLdE�vrU��[`�
�5�0��1q,`
]�^�D�i�Z�y)]7�^����2aX!*n�<�?��K�;�ZG&"�h��A����[��#�UA��\��J��PdU���Knf��37;��������S�.#	��{"^r�eOq�.�l�a����l²�t���A�)�Z2�So�2s1��Z�Y������o�~��Ѱ�++�-d�����Z����w�KW��@p��:��l��ɶZ�5J~Ǧ23X�g�iQ$��OHX<!�����(Ч�X_c��}8�8�Pj����}��� p�P�w���/x���o������NDGVK�wn��#���F)6�� M�*����@8m�ul�!�3�{���&�:�\��+F�˲t�Z�FŰ]������P6��Ĩ��4��$9o���t��٥ =�������-w�
��+��O"A�\ˡN���4�O��[����f0C�/���y��;��+�C�ŲX��&ʞ��H�V( #��bU��^��-�Yʛq�,q�� rq���bc��2�t�'B��T�y��	'ݟ�M1�7S���N��c�^�j��J��;;�氖:����*��/�tJ���Ų�p�^u�!�x�uYR��#��8=L#�g-�4��E�ʦ.;��G"c�]c������\�/�G�U�=�ܴۻE�4����;�r�HM2��[����zK X�����G'&�Zg�- ��-(��"�D&������4��0K�)vŇ{�&P+imvt�6�b����NG&����Κ�u����)�aьN-��Ƒ��31U��95_�@E�;��s�"���|'���1$���ۥ��6}�'�����uB��X��}��9g.%H]�S��"*<Ò�1O����w��pk�Y��1��w!r��C���k\A:�ڵ���p�S��,�r�1�@�?�e�܋�ӂ��'j�́����3��"[s�X ��p� v:Wu��� ����;
K� �������|��1�
��b�}��[��z==l��@wIK/a�%݀i�I�Bl�K�T���}-I	�1TU�cЭ&�RgO��� ̬Zzo!�y�M�߽U;��*vՑƭ�D�����giE�Y�i���4�b�Q�͛�F&t���b�]�/b�n�G��l2^�}��=Ά
����$O���'�.nd�^�: ��p�Ū��
��Iڷ���鰉�U����b8�^.��Z�&~M��E�ǀS�R��3[�������k��0D�k툾��T}仢S��	��s��Be��/r��.�
#���g^T#v�n�0J�+6�u4/=��Ŀ;�d�'��5���GD��h]��f��W�Њ�j5�WM�
�[@8��)��x���#+�A�G8��)U��u�`���p����͡��+n���w��C� �\]���V��ndc*1)*�S�}�Bd�ױ�w�<�M�G�e��K����q��ΰr����VU�����W볟x�@'���s-�5˗E�eu-fgq�)�~��*8��n�ŝ����@E�i'���m�9O"���K��[�6V�1�Yޮ�^	�>"��s"�������=h�FR����"�$���
���g)�y���#�>i��ӶU���Ѣx��9��w}��]6?]�r(\��O�YNT�d[��J���fBk0D;:g�o8t8�'�t}d߯�M��{��˙��,�*u��Yv�J�X4S�ųw/�����Aq�%��ߜ�I��e'̾?�6��;%�2�Q}�T��Cw�G ��Q$�,F����+���F�Ķ�z_�O z�e^���(�Ip��$}��E�^�3sGY�y��a=	� �qzƵ��E5j��ZL%Dj%���L]bv6�g�Z�g{�SߓlF}f&��/&[����C8�I��\�7�d�h���)�d�5��x�'O������#��Lz
hu�[=,���jv$tЙ����Z6S���Rm���MG�+!Xol����Lu��Մ�}�l�Xk8�m�O�h�U�Io��C]D�Fqo�ӼX�c��N��p /��I������XlxV64EB    fa00    23b0Q����'vMb��E�Ǩ��A�HYU�p���  "p�}L�Q����ڌ���T��ȟ��'~�,��%me[b�<ڜv��ZQ�hgXE�O�$2�7R񵺟g�j�9%kA�ΡP%�ōڰ�����Z̕i�Zv}]�߁X���b�X�&���¥>��hҴ5���e����m��y�t��rxt���p�~/����E�4O�z���i:T�18�E2t9��;��]>��Ny���y$R�W��E�=�p�=JF�v�`���/��N�C�f��q	A_����[�Ծ����­=��7�#U]?�^��ܼ>��pވes���̳����[��G�u��?2���)T��}q��i���A�Hq'�/��︾#<��"A�iD8�j,%$ȣ^�ҬK/W8f���h������ݒ�s��]�u���P����Y���W+)�[4�^�f����}�kptr��Ӕ�h滈�,%U�^�����{�����0rx9��v/wI<� 4qj2�]���Ku�K��'%g:H�3�:��V!e�_1�݋ȅ�R��DML��B���q����2Z	*�����?�� �����ma�'~�����&08f�q��\"�s�j"��(*i��߬tO\FOd��<�+[��KR�j'$���;����:dYS�1'<;4�Nzݬ���ºY��Z!f�.g��J�g��'6�0 �U3����Wl�~���΋}w+j|B�{++�\���mN�r a���j)đ�I2B0.�F�\^#��Q��Ŗ 9�!�\��Vp!6d�_���z�5O)� �^�"�W��,����{O�;6����O����ը��T��-zP�����,l����R����/�Q�ؐ�j�H�D��l�O;�Ӈ�C��#�`'?�K��&�]Z	Ĳ��i�2�j�Z{�{�ۍA��/>�9ev�n(��f��E�w7�v�b������a�\W�8�#$+��#�^�3��q
jy%;t��R�iݾ�2W��A	��_�xʘ��L����_5OMn���e3#iU������V�� ����#nA�}�$.}�Td���z�h��)��tC�����O���a��^�w�V]�:�ݦ5��+��[
�i�����A���I��i�2=����g㎄��색���� ��uPY+?��Opي�A�E�	�P��3�2�G^	��hf��v=�a&^��<Ex.��?�:߱��H�w9<j�b���z��Z�H�*#���E?��v��*Y��D;�C�l�= w��_A�����l-)-�����>�p�J�|�O(��[��u�َ�7���p�Ó����F(���Y	�DܻV����m��HgY�}�5��5B�����p�i���'&�߫P���d&��]�q���v!�[��oJD�m��Lk&�qV'=�m���$:&n�-�[B�TY����Z�W�s�yw	��eW�s�b��B���#g�)�^i��G���^ѣ3 �7G��u$06D:FFТtY�5m^��+�7�{U�8բSr�9��'��Vy�c��qr��ƪ���\g�7�g�NfZ���̍D�����.�k����+*�_�i,��E=C}B�ζE�Z�E_�����.� 0542�W�C����T��Ky"B�3���eb�l˭nF"���p[�0<8�����O�S]���V���kGˈ����q5���Xt�uB��$����P����f��qR�vi����쩱�Z�>��:�'.)� ɐ*��"睰��c��ŋ�"z�ڸ8��:d}�f��6�qM�h�W�����x�rm�F%��;��"�_�W�c�z�+C�Ai��V��!s!ՇB��.�O�6�!QG�-md1(��ኩ#b���cH��[7��	�>�H����m�vHJ�v7�x��'���oY<߅5�aE������l>am&#U���Q�Z�a:���m�*y����UW�oo�z�!mJ�T9��3��g��>�"��%bA�s蚶e�\�T��NQwf$tIA��%�UPf	�pT���8E$Ӧ��{���KR���	��5td2��P^ JsF�!�n{��!�o�MtW;��Պ���Ed����$��3�+d�{̖d�:�Iw��LoZ(Y���_;����Z��a%�7���Be=�������	u�Z����D��s��B	�%]0��g�uf�SA�
�|d�tz� 嶏�;B&-���O�+Υ�gTs�˲����q�R�Qȡ�K���-���$V�R���g;;�0kRc��RJs{���C�h�t�����NB���<U�L�H��}�OѤ�y�lTQ|z���Z0���'�4D6&��l>���C�؅��4y�Lu�j�g	-FOj&>����}
���� ϭ���*GX�bG�|���Y��'��������?$��?J<�l�[t9M����\�)�H6���4[y+��#�&�N+���,�BVe22	F����R���_��ב��G
2�.�I2�j���^�K��p�z��-��z!��� 7�R/�lK��*)����?��`C�|"[�E��!�B)n�yYU�weeFi����f��9�h���U��䴶��L{�@�I���kqb�#������;�ҍ�ud�a���ԛ�Z@�LJ̚~#��lG1�Vz�ĩ���<}$���}�A��8�)����B:J�ҶR%!}��y�UZ�r�h��zf��Yg�� �A�݀��M���B ����FN#v{��Vt��w~�2��ߢ3�3Ӟ�K����A_RS�ͨ���ș�x�;I"apdه��Du��$�K���]�0u ��,]J(ԊV�w�s7�	��9�(׮ߐx�0unI�3 �z�9��5���9��=^#���d^<�?�P�~�� �xJ�@*�� ����} Xr�����z7��P`oX}��p�<�FU].aH7�0zچCƝ%�����b�EB�`Z��m}�X�ެ?��?/y:r.���X.l�CR���\��p�VZ
��0Y��U�
&b�_F��@f���i6�R/��U���@U��8Y��\f\�9��*=��2�4I��9˃gD�<Q���i]��D�|o
���i�U�B���[uT�fG�u�#\Jo����0��p��h!���3I��d�L��EGZ$�l�Y�aaSN��qC
��$�  �	�sR�B��ޚ��AΛ�m�j*�7�y}V��YV`'3� ?�0AVjԀࣇ�����V�r��������h$������������mn�<�R�Gc�
���n!���- \3,���1]��KE+�"�MJtŎɊ�&�<t��י-���y/= �~�@{�E�u�_sT���͉b�3 ��rw���c�	ϛ"@jz����������<z�Z���y7+�!�a���|-G�Gy>�2Y~r��]��fhҜ�8P�"#�Q����N��P�͚q�ҧ�R
"�4I*�� .��5�����ʥ�'��K0y{mi(zA��/L��S*�����f�����U:��u��A s$.$��tW;������K>��Z�'��l�V��mo��v�����r{�fk�mk���.���Q޾�x\�v�	(�X?������A�e	p����{Ö9I�)��	_�KؑZ=�>�OT���4}r��ؘ�L�6��]_����p�ڽ��rl�K\*���ZCﳉxL�:��7�B�i���Kʫ��{V��3s�8$�5 ��.��߁>�N�tR��)?S��$p���T���_���WP+�ҋ���&�e(�ؓq��u��40��j2ֿ,$9Z���:d%�ȟy�8t�a'bi�WM�L�FU��5���t���@��C�/��V5���Rt�R7��3U����]��Mք����tlEu��xt����G3K��x�l�w,���=g��L��M�}��
��g�^p�2�u;���3 z�όk,�I
B/B�r�%֡�@_��[�;�<���,W$����5�l-��;s�#�Q6,�������M�!��8=Q�gi��;�ո�l�/���*�S�m)���e!��J^29Z��M���f|F�B�O^� �"��*�����w�a_C;%�&f�Jl<��;g}����Qj�4���ԗ#�j�!6E!�D��jЫ���zCJw"7���e�W�
�HVωo�f�� �t��/W��/�o���uX���
���rh½����v;j@�d]�I���:���-iTMYD��9��y��&�	���V�5�� �yL9Ȉ�Ao�Έ�oՇ@D(��Ht��8}xٳ��[L�UQ�y��^�B4ҳk���*��N�RJ���A���~n�!��1�>��ɰ�[-��<,��N;�`�B��
Y���y5>�O���'ǨC�o0��H�ڥZ>p$�5C��"�����Xv�,���f�,��bh����l�f�}�(�li9'��A�Q�Ie!t�+�Q���&�;�����E�³I
��dx~�(N濓�w�+��Pd䀋��XM\�}�y�a�!�B����~�(�ۖ�_.nB�Fs ���A�A��y7S�(3������Z��A�s�9�����F��hj�
}C�/���7����o��pj\%��,�>gɕR� �?��	�7��焑;�\t�y��х���f4�x� ��\����dH��d��~���ʳӛ>�Z��v��D�!���B���q���g;aT��g<�뒅7��QD��bdޢ�}0�$��/�f���)���i0hޡm괗��&A?��f���z�T�p�e�B�	��͝d�}u�Q�x����-�\^H�Ǌ���8�nH*��n?{�i�{EH52�����1z��P�(���H��d�BbÜ��1�lI�j��Ҹ��Pѵ����z|��ԋ:����lZ��M&���d�aM�._y�R�a�`����ZfP>E�[��d�m��f��DT�Q�_����W�R�����8�d�ǻ5Sq�}W<���O/Z�L� �	1ü:�w�zPT��K�Z���t">9�JI�:��Hdp���� ����Y��!�	������P��^,�<y���aw��W�t�˶�� ����u���;�.]�;���6܂ח T�{h
=�#�ئ5Qqn4�&q���h�pI����3��o�-j�"�l�Xna%� I>|���
�ӥI����|�%bM��WNsb��D�#q�Co�AS?`틜Q�j0)��8v����Vm��#j2z?�a����y���FH���Ng@	$��a�IH�t&r�����m�E�_u�5�}�YC����ԣ��B��7�#\���c����9ϵ�5�a�ĳ�}��Mf����gz�����=8�s�s�BAݷć��0ć{<��̊a,f��U�b�����ҽ��K�_�l!D�;�GL���h����ˁ�����px��W��7�-2n{�e�`��U��A0��].+K��OlK2�g��N��^l|
mf�&�0ڗWB}��|�	t `^XS����|r�f��s��,z���j��t�5>�ӂ����e�k�tS����3[,jO!
O�j������@9=�i��7p��)k4)����u���$�F���YMg���̀���urqz36���X����b8�D�P����C�	��_���2;S�zԵvy���c�L��`�iKD~��Jğ���B*Q�N�U�ޝT,���Fg?������f�UA��UUJm]�ـ7s~�xa�2�� �>pyF��w��On��v�pE�ņ��5�5(Թ3����}��Lu�'z�7������c��>�3\��t�����<���7�Lݰ�&v��Ԛ� �a�~���(Aݗ�ǧ!"�c���8,�ة��?ζ3<�>�ӄU��z��`D�!���2�/A���F5F��R�L�XS�A`}�^0|yeEߌR���\N۞��j�Nɚ4(U{��HL����;����t&��e��� fjVQ���Z(�@�A6���%���?�=7~�F�D�dK1A~���7ē&�9�����n\��|�TN�y#M��R�5���zT#$�o4!���V*�x�E���"+��"A�\�~o��r��4�|��E�?���ܼ��g�[�z3W��ߘ��s�������M]ɪǨL�P���rk�-����?�,��ڮ$9�2�>m�|L
���],��. ����x��R(�<��<مݩ�=�����[��΃H�ʤH���h9�-�{�����UI\�a �"~0?�冒���v�� ��\"��Qr��y�]��>`W�g,�{�Z�C>�����Jmz���yp����%ia7�t�(<�������)ʂ�ȗPO�q��F�S��X�%\��d��lt����d|�T���ɝ*L�CB��f\��@ѱŦx���D�k4�/+��\N�[�N����Hk��UEz��>�s�w�炰P��c0`��t�G+gi��٪�[��b��B��e�yMD��LEC'_�"�̇���p���YUd�Q�||Q����[7��l� �N��}`t��Ֆ���p߰-
f��v�Ƥ $����*@H���l���}����k�0E�>F��M-3��s����� ����Z��p��Ni35�$�`TN�/��3>Y=гB�6�A_��CGE:N��C�G�S��z3U�=��t�U��8k�5ZԦ����YΧ���o�Fe!X��3�$0E�˦� �N��u�Y�P�T�x��C�6w�F���%k~0��^�x��=� �|2�0���"i�Q+`X"3���3��9L\ݕ��#�u�<��5e@	R��o��T�炎�Y��/~Q��f���தu�_dp���׀�Z�XZ���ַsV2�܅$h��<��kN�UqW��{$�A��=]����@�}y�5��D�Q��l�Lv��vP���3jt���;$�6�O�S����v����6����Z�>R�g�aP1m_B3 ��@w�\|�ٴPq�~�T���M� ��\"���L�??n���}0}S]�q�B>;��93myB}���;y���汑���d�,���u��3+�d�e��{��XD�MgxFR��.Hc�qC�%;�	 �h�սKłg&|զdE��~����>H�,�K8Ca��|_��.٨���q'�j:��622F$�	�\T&�Zѿ)Wde�����$SV6-�~�wn+� ay�N��I��R�4|���(HA��h���M���H5�����Gڨ:���{d5�V&<����ۏ����	��  ��B����Bf�%TƹCn;��yO5�y0�� 8�Et��4O�ut 7#�|%�/GOF�v�T4��܄�H�r��D�ќ[�����g�E�H�\�&�����m�A ��s���k������W1ŉ�����%�����݊)��aND-I���q�W*H� x+�E�u�2�OS��6�x�+�C~�a�q��D��GPO����UgJ'�h��u�$a:�m���;��(�ѡ�&#��xL�&,;�n�����e��h�� ��uQ
�Y��I?0���.   шa��=B󵔶\�_��6C|�&��}�0�>.޴�f�|F��Mk>푆�Z�B���b�;��99/�ט�%��x��:2���N�ט������!��k\�eѓ%��u�-0"��<LW�0&�������g���Uv����^
kL	�cj�v�9$C*K"I��r֏�7�J���R$�3����G�]c��r��-��7>`���*�9���ٟ ���!b����oݢ��mO�q	E�yYUT��d�~	���k|��� 1��d��>+����Sj
	C�"~8���bK���j��T��/9���������b�Ng�$���?�6��wd�F��������X�A��(0�,eB�A�H2�*��!5�m)����y����K���+�Z���[F'EQ��.[����?���F�'#�_k�z�����#��!ʒ^V�Z[�{]�LD=��b*�,��������>R��, �Rnh����^����Q��
}\�N�eD�/�<��/e1^dcЃO�g��K��M�/V(�y ]ݾa��$�2|Pb�!��K�d�<�b���Ļ���l�_b;��a2�UK�O��	�\b�`"�?yХ��vp��ί:Vc^��X�+'���G׌g&�ZZ�0d�a��䋇���`1��ў�� �zneDj�2JjrR^9�Th��#����%�I��&�5V��Blt�hnY�JL��w������[�E��R�sS�1T�=�����
�k.��Qwc�aLhI0K+M��<ˆ�35���C�c�W&���t.srt��*<�7���n�㎩t8�w�/5#�6ޝ������7-8m�tB�ı�EWBi<�
֍Ѩ���i�gS~��!X��0���ĸ�f�C���#*pXiJ�������8�H�[_���=c�{fh4����GAc��8Ls��i1�����d��7�m�"3T�o%��v-��hH8�=t���A�G&��ڸ���0���ڟ8Kd{��|�01�Ⱦ+�ek�M�L��[:'x���ô��p�L�P�uOP�c�v��!�gI?
A��bb���eI2�/�v$D��(��q�c�d؀X$��5����������=�ܷ~߉o�1~�*���f<W�ʙ'x��[J0���+� ~��h��ᥟ/oW�9�:xALw���S�j.}E	�:�L��>�+�m0%���pWf��'r	] KL�U� <��\^%��g�%��!���� B=Q�S+�����`gЊ�{O� �B�����D���f�a��0|Y�!��T��i��Tb��!`>P `��̄�e2�8P\�ύv�j���=t9�����S.o)^�9?0��^�� �-�y����A�c�5��|!�"`\���(��&UXlxV64EB     a1e     2c0=ԓ	䏎����m��m����Z��s�o�fy:R]2��S+ڏ�_�K�Ich��(ve�QgW�rU[�׈�ܹ\��h���[l1����q����G��y�ϐ�vS�f�We����#~�J�zOR���&ċ�.~Ug?��n/آ�eMG�j�_t4�
<���y��n�z���et-T�}l)������uZBX���X�剏�?�Xƌ i�^�3��Ŷǐ1o�X����҃���+�ݡ��E�Q.70U4Hls��.�eE =�5o3��	ô}���<E	&���c�<�n���q��u�J،J\�T9�9?r'�^�/c�6*+���x#������Oc�Q�J�7c1��2���b�T|�[���
{R9�����*O԰<6v���'ߥ�˴E�:l<��P\�4' �DF{"j��i���U�+��̔�}�~�g� so���0�l|?RpY����6�~�l0?�!��ng�˛�|O&�{�m����3tG�Z�w�Md;x�x)b'�S���sm�-Q�ap�w1�_��S�^�Pqq�,���=Y��^n��}(J�����-t"}�����ŜEݻ�`��'������Op�n��!=�,<_!k�5��+�`v�)�+p�E��hp�����BE8�1CT��g=8h
���K��FK����51!,�(=2)%�