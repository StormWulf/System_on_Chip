XlxV64EB    25d6     bd0h�_8�b�X�Ci��4s�X zv޷LX�[�M'�����c���.�F�L��֥�Υ��f����Q_�T}Y9hL攚�b�	�#	9Yv�9�8r�VhK�!X���>-�e�5xS�v�ǀ��X�x��5ycrC?u�_e���L)��+��i*���qT���>��:Z�~��{�Ӈ�<����m� �����,�>����Ъ(Î�/#�y����N�#��܌�]��wxJ-\�i֟�w&���]�����ڬ$j����~��j%$���[�Y.7�� ���(?6I,"�O��I�B�
v^��a����D}@�ٻެ5P9�̓ J�1�mUA���Y�Ng��/^��LJr�d'�V0�@ k��,���Ye����d�VE;G8d/�^L*Y��
g����P�C��(�XP�2�n����cB0�q��b(D��M�ͳ�n��
��W]2^���Ђm��k%~4��m�2&1B���dD�y��n{��F�I%W�Ƒ7��Ȯ�Q��5�������P��g AR8:ѹ�����6x�����4X�esfH���α��lv�po�NLj����B�7�ۏ�~j`���Ȩ)S:��Sh
�S�.�p�x\���9�)
�f�vi�<ً�K���y���(� cHp���X�@��9+1�b��wH��q�Q7 �ʩk��5�J��  ;w`8�S	8���A��CzB����]b��z9�ʱȪ/+���2"�6Ϡ�A���J?(���eƄ�fN�Ւ6�Q��D��]��܇�y���*CS&v�2l��t�ȿ	6M�%yw.\������y�4[���[	��p[��<ׂ�mo����R�P���<���.�_~�'������qKN�1�ǚY���oVfy܁V�K���o�O-1�Q�hHz#)z�k]N���6��=/$��Z뵮��rӖ�u4�R��Ex�)��{�X�E�n��~�H�^�q��5�B�(����bӑ%f��/��	!jF��_F3��������t��z�B�< �\(j�]\��<�[qQ�������|t0�,Q��낾N��+��H½�Bv����(��̌�����_�S�������u��@�����>:�;ޡ�ŝ�7���L�qs>��P��e�h��I��7(��40�f����`�_#���*P=Y���نj����2�Z��s��ђ<<*�B��G��kE�BZ�۽%�}w��Q��tm(�(i���O�e/����� �<pG�7�e{(�B(��V�����[�o�w۔��ܦy�Ρd����#�vc���pw3�3��+Y���Xex3���gw�~�ֲ:nt��s�f�9�$��f�ȋʹh�C�eR�/���W�ҷ�߲�A���]�o��\g��.�&������{�6��("5�/Z�� ^�h�#��;^|iL1��	nc=��z(<�xK��Iu�ÓnG��9��0��uF�,�5�H�Þ��a������۝wI�3�H-�{;|T#��h�
�7�PKk�n��GuV�-.�c�f��%�So��V��*���3������2�	����5A��`ϲY/Qr�z6�ۈ��� :�^[�L�������*�k�2z����-'�S2-��߷T1r�i4&�`�y8��]ʵ��s�Vc*�茁(�EE�$���7믌]; W��>�גGa|�t =V��HO�g������6����wV-������HIӦb^�P��Q�ͺ�!�Y]㺰~�[��@�Јް��5����	��&)�����5�P=c��<�	 d>�>n�����b>M��#$��+] ���S����w��1y��v"��Ƀ��g۽���!2v����X]>����3'�tK9�%��ٸ��|>"����ˀS��V�h���cUT�`����vj�=�S������f�[�Yt�"r��4�;LϾ�����
�m)%W#�c�g;\��b����p��5Ţm����l�|'�LX�kܷ�����]�]����Z���c�x�_�����p���������`��D�����y��U@I�'����`_;�"�2�C�@"5��H��!���pK�C�n�]WY8(ْ��>x^y�W��{���%�D�	�n'����=�刅7Ax�WR��4��S�6�61n�`wM��Uؾ�ӟeҋ��R�,��Ef6%�l%"S��<��Z9g�z��d'��XA�ٯD	8�d�h\����/���4IcADעE��1��v) �&`�Gp�〞o>o[�{mKh�!߷��y�k`�+�]z�[�S��}���7��6�K�Z>�'$r�*U�F��S.,'5̘z����#f�}Ba����8�K��XO�����U�2���K1	���>�z��_��Z� �
x:���N��`g �$�qbbgI��˓2AĠ��-`�z��l��_�j��qjbR�A�A����%\<�l��GR_��Kr�N �퐥��e��f~\��8���u�8ĳ�w���v�$��~+�L��3�t�:N�;��D�ߌ ��DP���Ԥ���������H�a�XЕr8���^(�*���4~n���V�WCY�R~)V�e��������N������d�;�.]j�_��3�_�R�Vj���5���#û�C�4EWܽo�E�'�"I>;�KU��#)&M�#J.����H��v�<�	�&�==cRTPP5�I��&a�AB����F�w��P1�y������"k-����f�yr�	ղ��g�9�P�F|ւo��^(?�������T�ɽ3m�in�E����2��&b� E6%��9IO�$F9��ӣ:�o_gAѯ˘u-N��� mth� j[C��Yd<Q�3����(�C-��v�PM5!��?�t�#�,@F�[4&�Xp�"���b��{7�R*+4�"��f\���B�޸JP�p��Z�mf�H��r�FV�������