XlxV64EB    576a    1430��Z[�v����h0.B����{7 �vo�]�F�S����`>x��8�C�
��Ⱥ����� �2y$���<K{b4`X�������bԱ=��}*!�J9�[# �������SԦi��r\,�`0�	�g��]Ɵ6V�)��v���
D�P".=�p�<)D�)\���Ve;@�&��9�Ֆ�iH^��}��L4�����RUTmS9�8h��m��q[a�nVx�+-�z�(�=�<9l�E� �\�'��G�ɘ:���9x|y��z$X�0��(.0�캻�l�PVf'{q�*f�Ѥ�p�c����� W5��R�����u�R�^��t�hq�ʠ��"PEqb�@��:l�r��'�sSW�3I�VhH��#�I�q��".�j�	$�|��@�2<�ںbdҏEQ������`M
��=4>���lT��A��3�M?��G�cM��+���P'��IM[�����Z	p���E�J���#Zz���pQ[i�F�{�<ۯw��%UR��ލ\d@�+���_������u?���s�U����Ȣ�CNu�z�+�zcg*���K������@��e'P��Wx�3ֿOg�d�F���)	R6��ֵ[�dB�v}��������Ɩj\��&]�	D�=/0]����@ti9�Gd	�Be���oG�Q���(�v*|�@�j��#�jIjn\d���y!�diT�g�̥���+�G�$a�(��������Z;��x��:��3�={6[8*��������N.=V���D-�;޿�js�:|��A��\��؝Fe��<�7�5���gOx�>�xnY��˴xF�L
�y��/�,���K7�^|� �!�}���QbA�i�-�+�������Uj��t,I��2�PɎ�=Y#�5%�KHt��0�����#U��/�� 1��ܾ�\OϦ� ��y��ws@�P�8qy��������)�o�~"OB�~�I����F��N����3��O�wT��(#t��^�';o=����}hY�X�xy���*�C���7�[��vB��+x:ݰ�\���Օ�;�i���i�3���`X+̓F�"��5��L��V�;Xa�7nGs����w�:W�Q��0��h̹7����F�~���Ӟp�-���$�+��$�ph������$�X\�f����}�
F�E��@�kЖI��&ӡ>��D����/]�1U���튔�8���I�?A�؍��Ն�f)��!���z�2;1�� b�j�|x���/N�R3�����wJ�������mځE��?� B6��4�mu"�f�F�N�#m���/�5+J�V�Ph��`fg���r	�W���Si��tɹ����}�"�8Sc���O?�םy�k"
1^���~��^������,d����/� ���J���� �g�r��\q�F58���u�x��{Cgf#Q����K�����LG×���C!��x�eH������_���-*�v��bp�;�Z�iz��nM��Qz�Ϊf�a����ZL�.ׅ�?�o�蟯*xt��VL�0r*� br�g��m\"����b�.��Z�I9&��j.��z1�Wꃈm�d���<�B�b״Ў�����/�`0x�3|z+�eP%�ĠD0j5c�曪=�K��ZrJlzyeG̤6�^���7�:���	�c��&x�ö�ڀ=r�;����~QN�c�{_J�Z�.u�ax��5��eCM�o�f��p�)��g�ap?��4�D$_`1���<�w�E�3J�(��l���������;�%C~�'L�_B���I���kU��2����/7km�<!�!���"�K@z��G5���5��G��=���؅,hoL��α7)�%Z���N�j.��t5:�)�Κ���A������zb�5�1sR{��%�[)N7"AT�������y��<�h�q>�_�{�n�� �\c.�͆����qM4е;od������(J��:)����ڋ䙝,Xj�Ω�)y��f�g_Bz�S��M{}P�K��=�&�3�5� ��}&��?d<�BwW��&`��A8��_;%\P�[��\�Qѕ�t:@[_�!����:x�����2��v��[V���9��'^r����_��<��[�+�!�X<��OT(���ޱ�k&6�(�&�mN�|g��O	~޾7������`L����d��=C��p
]�51!���Z��<8!��P�.D�8���15�����Լg8j�k���2��~��|��p�Yв��bD��jW�������k���$r��R�e��E�����a�S�386��L�~�u<0�u�)��./LQ�� /�|6DJw9EK�9e5աw��u���7~M#�w!M��ˣ+���ɐ?ӗ���AY�y`޶�u��=X��T]��-j���m6��ow�z�� uv�Z޸��0��\����)���{u���>Y��y��
���m�йh��{��O�e��+i��Xf�tǙ�|n���oe�7�W�f�_-=��P��� a����P��ZA³��+�#�y���{�g8!f���,㐨&rQc��VY��2PyZ���qeCj0C�,�w������X����,�j���SU``y�4�働UvSl��3��p��=�jiX"�<Z�`4k��k����2Q�\_��#�4T�܇\0�C�i���y�U�ȅy�.���^�d?��:ð%&�J���R(�[��!^
���Zm�4դ�ga4-xWK�����Q��� �ú't���E%�K4Y��p~ϔ��hz�'�^MN)U�w�Z$؏��=R��H��\��r������bDIq�&1�߈(�� ��pi�G��0�����?]���j����zY�1�|�:�A��o��M���5�^��#��q$
�d,�ѥ��%.��>9���=��z�O�F�ڽ����T\
f��oVE6f���f�Y��T��M���y�
#�Z��.���<����`ocs���&�<Sa�ŰhXE�|&�SZZ߾���'�팤sF\4�:Lt�R�6)l'�*gְ)�a���籁��]���~v�����>9L��$�@��i�v$7R8���%y΢=q(�����1�Ӹ�d�%����-K��&��#���^m����"��Ĭ���r֬ow�A+�ʂ<�ۣQ��m� �7"^�]CPe`O6�����7&�q���3�5^�+OpA�ƨ�^W�v-��6ә,�E��(�@����z���,��L��9cAVL���L�?̞�1�<FBo��ܬ�܎�[,'���
0Ȑ��4�
&HC����T8�.�����7w���e[ݵl�ntm	��"���
]��	�����R֦�|'�����q4uVz�Ф�Ǐ�`�26�?9�`�f�`э2tn^
&�	�S�si�1�6��m�@�.���6�
�1/ߊl]J�`L�^�H�%m�6�Ï�8űMݠ��J�dJlX�j|��g#�������
��oU��W�X��nE��.|���et^7۟���c�j�9^�E�B��GU���*Q;�^��}Lk5||��~e^BE���P��B�C<�����9&`�i�����KFn�qd����o�W*O^�PDq��-�T��%����!���QH�I�7��0���P����Gg�ĺ@��Q�*�+��o�<���	�����HGB��K�q����u��@V*�ɸ�;�zh������:��o�-{i%$�R��R�}G��r����H��CJ�1S��9�<<t�x�Q�T�:o��a�ߢ�H�IQ؍�#��JZ�J�:F*T�GU/�KiU�
��lQ٠YV�3�p��v�(OڕEf��wN���#�����h��+����4��c���.�͔3����� �cۙ �RvL�e	�t����z�Oe�c#�����߀AAz�T��~M4iL��Kć���efQ��p7��d�	��~qv�[�W�N�DNjȎ��E�T3n3w�չv->V�{$�>��~�fQ�o�Q���҇P���X�N{�>GJt�w����@����d����F���w���S���'F����5Y�_�:��8Ko{2hyX��\쟶��Zb�.��?m��(�n�(�-��_~�W�P��k�1��M��\m�#���<��r*��=�R��!�I��79B�%�90Ew �}�|������6�UN�wu��W!���Q�,�W��La?��Ł�6Y�Gƾ�6�}ӅS�诹�W�sU�1�}V
�Q���-W�R:\�*�\��v��~�r�9���v����/�=�B��-mQ�$d[�fK Ǔ��\poJQ�=��JK��
�b��V�II��Īd�bF^꙱]3��VR`9�:�R !�*v��Y��w�v��x^L��)Kp��t�^f�=,n9X��+�z>�T^����ፊ��E&{���[)��<�S��j�a�P���� /*=qk[���|�T��͚�]Ԋujɒ럼6��@�u<�b}�f��m�jTY����^�h��lb����g���9�#8FZL�E��n�&(~�|����F�s�+�T�5d�/!�=���_K�K�i3v���<Q�N+���Xa��r���5ƍ��͇:(�I�*�5�laI=E̠Q�(+Hz�P��2U�3��^��N�a�$%�#˗�L9zSbc�S�t�����$�����Q�g�Kā0���	��*�\�P�S�`���(���k�H�F�=�m%���x���D��fQpֿLDT�}�G sGj�?'>SK��c%r8�+!������c����uY�JӚ��/s��7��1{Ր�PW�m����|zY.)���X\vv:���n�8Yɖ�k���4�La��C\����;!+��4;;�`��ds<�T��sAާ����|"�"���k�?��yG_)1�K&���ҮbϮ'�b@n��p:0�/lv�d�WΎ��wQj	Csf���{5�Y�Ǿ�U��O^#�b�TB�覆��Jק'�A{��_�E5ʁ�r�W��2��V�SQMD�]�3n�M�W��R����Q�F��XP��C�	���Ofռ`�js�D�f���z