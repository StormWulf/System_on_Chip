XlxV64EB    820a    1460C��+c��̝'/<S���J{���H��8�`2>��d�B����TS[}$�=��QHUB-�c%!Z[�D(����6�J�G��;^ ���%�-�� ��g9�\��E�tٛ�O6��`���e���F�
��V3߭���g��{79�����w���ßuM(���	�r����d���|��:����`w}�Ռ��S�	L�2JL�{N�{G/��
H(�T HS[���t�c�Y>��X�TL(�\y]�m�٩ڵu����6@;b�s?����j��P������kψ	���VPsQgD8#���j��Oo::5��jj��s��� ��5>T���BO+�w��4�Xl�}�:�+R���6R��'H��|���Ui�n�O�d����r*I�D{\�[��5��d�v'��4�]wi�b:��u5v���<����d�bc\��=�Թ�����̛�hWn�.��|�n#��g�|���3�t�$�'�(�`7���#��gb��Z���+�'�=�:$�.<�"_�n�Y�����<3�j,�S���0�ֆ
e�]���'�Y��]
c&eq��Ję�/��;����G�O�����;d��UF�δp��P���Ĵ�%�K�x��"�I�@��u��O�����'�uZ�!�y����#IuDRO�4U��߫�d0e�̋p�����3����DZ<lC5�*�R�S���W[K�FG�N_����R0<���_�ͣ⭆��_�bqEK�����-D����(pHV4��qHu�����R�A�}�7e�����ɹ}]�p���0m�L���� �nԭ�C���2P�b�&�{� 6�Uh��R�a�#�� M4|9�hפXs��K�B~��⦦��W�,�)�H(�$d'�N�J^���T��ɲ�gj��[x�m��u�6�n�u���\�h���&+�؏��(�����gTV��H�v?|�n�r��ɶ�: dC׼����4b���A ��6u�]Nq�5�꘭�n^�l�;��}Np��J����
���U��~�U��!wZ��V��d�"H|/Mu�Y�O�ΞԤ��E#`;�V�&��� "՛�-N]���/lDXd=�{�$M�+��9Y���h3���L���h�b>Όwu^d .Pa�N��99V˘���Du0U�N%xH����4|m��M��۞=dH#�="������u�L̨��Y�dW"ٯH|6\{��t\��߉�|�hd���­l(���j����!Q�{��-^.=YZw��K�zj���!����U��(ё�I�GR{J4A#�aʸ����T���L#�b��+M��:��]}�຺v!z�K�F����&�������1Ե�Y$�F%f�On7
���@3�S%"Kb0㵪,�c*�Zl��i~4��� -��#<�N��'�RBV�Z�Sr��hS/�F&ȁa��V��6�-�3������a5d�ŹjD!�:�]�t�̏x%	nJ[D��9��׌`/�p�X7d�$F%��|�.S�������Jٌ�"�-�����V7FV��:]��)��k�` w�x�=�j���LMVbp��mG�*N -���f�$�4�y�r��SI��e��\���{��Դu�/�1��ʒ����y[��G&��|���]~L��N	��]"��4��=R�5��s���:��=�,���Ѝ&�<d�����"H�;oa�ξ\�6��J�A�=�5f{��=�������kz����=���fHժ�P'�C�陓Cz���^dT͕
4"j���>�9��F�ѽ2o�"�g�F�٣o`�?/ʰQ��@"�`����ܽ܌�.��C��ly�]v��7�	��'F��@�r�r�<�\����>�w �1�ͫ6�}#�&b��Lgg�-�]-�����������z�e�����w��Yp�Dt��$�`�̦)tov��~� &?t�)}ye�1xNZ(R��y�*Z(�ģr�S��$1<Q���R�)���%���дp�^�7���^"�=4�uU������,���Ctp�D30���t�@Y���T�-w��v�p� �EI�f�_rnB���m�'��Z��$�q�S{+��c��f�	�%����10�� I�8����^���X�]�?�+vE��x@db�~�"9�L���S7*�utO|zp�!���Vc�]S^� ����蒸�nD`}�����e�^HHP8LF�ǈ��6�B�%N�{̃�@�6;J�LlIi���c��YS�
j�xTP�\�P��C�D��8X�6�D'@�ח;X�pb�q�xlnT'��c�7#9�m���H6���e77L����sܹY>�Ԝ�(�Ie<���aɆ�.`�?�-]���� ' W�]����j����7�w�Wl��w�<S���ETt=��.�$�v-�	��1#?���E��nz _��|\Y��'��м��&�t����HQș���X�^?���=�~坨$��ƈ7A8` ǯ˅>p�V>G�~դu�~~�E7	�S]��R"��Y�5'�'��(y���in��笶��t�A�tB�p�<��J�VC��#���O��e5��+����F�Q�9�H�E���X�L��P��w�(�Xp��
h��>���Î�d�r� �G��A����f�4}d�k�%���)�%���m�v����0bO�.��#�
���ϲ"�\}���~���e!�0�� �;�o���������T���5Ƿ��Lk�O��δkA�t
��ͥ0^<��p����7�D#�Ͳ���0�H�*�o"�Xγ]C��!���!�*5j���(�ɉ^����m�>N�
N����bB��ME@Ny�2�j9��Ԉo?fa��9X�*T ��s�W��*�3s=��Dt|�>?zXS�R�$�zx#�g�VF�u�֐q��\@�km����m�U�f����*��xq��GnZ�XM�!��v��������ؽ����`@��Q%N�j�L�!�V⦋P E�.�g�[$ �]��	$d�Z6.��}r~3�|�b?�}a�Jv��6�AĝN,8�`� 6=�Q�bP����
��誸0�V[�h;}NI�D��"Ts�I9�o�zp����g�j�𫼧^��y���f�ݩъ[��j?�NƱ\���]�mEb�De�و8�#:NJD�V5�sd망��I~�ɛT�cBHfH7��[��%����G�n�R�����쭕��đ�I�s[�W˜����,)}j<J����h��/�~f���a���:7mev��v���GΝ(s���}8�6۵vNm��G{rH�#�B�hʹ��]'��F�0)�'M< w�D�ZhA
1�P?�~3���Ñ��2n��׸}eA���ot��Ӵ��ha{�Ue5��<�d5�r�Ԭ�w
w��C�֒��ʇ{J
��D�`�@�����,�w��)5�������{e�ｚe�^!�����b���v 2���t�qV�<���Ě����%��[j���a�9[#����E� �h*Æ=Ŀo�N���l~�<_��Q�_f�������-="ѝ��1�V2�+V�W%���om�f@+z���H:S���4D<�o��+��?=�0>Աt~P����s���o<�)j7��&��q���Ҙ�w�����j!��UE`�f�ŋ-� J��D�0B��Vjbٞ�;=��r�&�|�L\(���B|T�����򫲬v>�wtjٕ��on6�U8?+��{N~�]0�L�5���kc����{�wۓ(�β��Ͷ8q�z���K˸�@����^,�;��G�cMq�Xh]|�v�>��8�3%���E?AdvZP�,g$��<�)�JL�g�(��^����#F��{|�kÞ�7Y0�'up�`�(�1]L�J�<�R�V��-T[[ҩ��|q�èi�rs���$$�ά.�_;S`�	s�T��R��<��~Tϱ���=�����H�cT�8n�byդ�)I՚�_Q���{k�h���F��+�����|����וTJD�O�N�,��a+9������!�X_�30*gRؚIe�����a�$�w9l��e�h�8�קv�r�!A>"+1.�/uS�O׾��AEp��з��`�P`g��e��f2����9�%ض� ܻ��M�G%ЖN�aV,�$�����^���V�܇��+%�A#��F�ӽAY���2-�Ñ&��kE���}x�J�b\��1{���P!LP��3g��w�y�d�N�
;Dw3�a�_�C=�\�	j��|+��`�
z����Ë㰈�S6�8��qU��p$�g�X�t�x��q^�f��J��"��?�l"Þ�ݫ$�q�y/��I&�V�l4�:�d�fEP^	�糼���Y��o<W�?L�A�r�����^u��Mc��qYAqbS;]W4LZ��S���6'��St���H�v���cq��܅͢UR��v""�=�$�rV����8��"4�_���Y=;ۂ�4��h.�"g7/ѿ!텵8�Ĉ-/�L����k�:S��/N?�goA%�Ӹ0]k�� ����QC�GNMm/�ۤ=u�aLf��sB|��B&T���!�3���.�����^�}�	��Hk�=����$���li���&�������;�� ����>��"�O�+Î1[}G��H��H�^ɼB18�\W�qIC��}�
�t}��t
oM�I/�?m�Vc��sB:?g���n}�ȩz���n~�m5I�,x���Q��]D��8�Ɲ�a������7�ta$�S=�{�+}�����oY vhMG��h�P�M����P8�A�-7M
�����u-N�o䦗q)w��M�����- ������>�/,�FH<��Ԩ:�	���~�'�^4&kn��y�5�	#V�ƽ�Z����,���6B��*ZGH��Sx�a�W��5:�Ѐ�]'-&��)DǤFk��<�@�R��҉YKB�S!ӿ����s���R���c����J�ȃ}�)Ja��f��&�[q��~%�uP_�3��mטt��߷/hh�^��?�i�n��`�^��K:�U�5q�Qa��?�ō��'��p�aߍ ��¨��]�"C�E���%��[-� 0��F�~�N��<��0�Jۇv�e$=���x���`֑���