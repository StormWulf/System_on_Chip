XlxV64EB    2e73     cc0��8PQ!�Ɉ�>�o*�'g�d]�r� /�	$v������W��4>�6����)q&��R�$�ʜ�������m���1����~�����Zq���������#�\Yǂ9z�|(1�޾<�lj��v�"�O����fS2z��E�Z�}�æK]���/����F�K�k�����ϹZ�(���q���\3�`�=�;xK\��G[$6�xc?�[����^�ӆ��q�QZ0|@4�7��/BJIV[���}ƛ�nD���M�dӻ�^mG����K=2�N~, ����};?ھr{��,&��W�P�Ǯ8�=�%�<��L��EK�0R�C��S�Rz<�ˢ�|��'0���Ee���Z�(�7��y]�D܅�5���^�U^�*J���Z0/�cd�`��VeD-�x%�Y� `���ԩ8�)��ߞB�;��g�t#�ZxJu{�5%1�Ps�$�oT����E�_�y+ܞ� M!ᤉ������h�GC��w�T���������d�ư��
��׍�����?p* \�h�g��-���b���(�'�Գk�0�F�S�·�^=h�@�t� Q���Ax�.*�C� �tq�mL�o䧗:E���J��dm��Q�I�b�	��2<f�-F�ĭiS�+���.|�)��_Q�*t^�0���J	��(	�x\'~{�>y��Sd��̶ �DGv�]��|�d�� .�y�ٜ*����
��I]�!W4j��?�d�N�t��8�1@L�*��c� ���D�k��ŧ����;��!�5myШ���H2�ϡX@��VߊLL����ې���G�»��Q�y�F=���z����1A@7S�B�c�w�]�y�.�Vm����L����ř�s�N�0�)��Z��O�n����/���)O�����f���q��s��j�hDH�N��[��V=d��u\��(����N�?Ч���ݶ9`˚�Ȓ���c�M��?�p|H<��f;�>�A�;�&ky!?���X�S"�!���$X4��P����ܠh�˳1�efR�rjmڤ�)l��9�.bGfuB}�(����l��a�N��^�J��͑ή%�v����i�^�M�A�0�M�f_M�TƏ��ohRdh���H~��5J�{k�k��N�Le�}���r��������ݔ8n���P�����q��	to#��Y����ܱRu��!��R!��v!y�뜠L��9��vwLR��L	B##�t<)�gʊI刕w��#�\G)�A����cұ2���������a\^�D~�����\�h��ł0�ݹ0i�N���_���P�0;�֙Ԥ�ye���PvLO��Q<�)E�{�$Da����ox����ٯ�\|�v� ���!��Z�t��_�R����\�ił��V��hǋua��]h������Yʁ��o���>ዛ�'�)��%4�(�
^�oY��y��;�A!�:�Mp��V����r��ނ`Z���aR�b�e��`ؚD���e	�޳�>���E������C�n��:v6�oy�����e}П/�d�.!g�Jj�DZP�&T�#��-o����p���@�o-��r�w;�O�H�^$>��<P�Nx�DD����+ ��M�+�͹�(!L�,����Kwdv�*�ʷ����N�Ł�\���N�=M�_�����<������#ڎb�P�*% !��wBc��Yv�n(t	?������T�4��4"Y֡�$�,������Ua`�ǆ:B`��I�P�T�Ck���Q����m���EkS�T|�Cd�)k�(Z�o�8݁�J�h���p�h����ͯ�s-aP���2mT�3���N4�n�Ŷ�υ�����a �G[C�[r�y���x�)�	�v[�L9�Y矾�gϫT1��^�8O,_��APn�5�^?��*�3�蠹�L�'�>�ذ]�ؑJFhj_jѠs�Li�Z�ڂ�A�׍'�.p�ʏ���!߿mBt��G��x��G\���@�쥓jV����ԍ��n��0piYP�(���ڹ�͝��Ms�b����u�h�%��i�v���4�)LnJ~��)�Q�3I6sIQ���4�S�[��m0�w���4�6DjH�UrA5��bE�T�����Ԕ���Hȃ����2j6w�����o%�pz�
"O�~����ß����9��`92
{�Yl��ϔ\w
C$���[�%����VM�c�a��h����݇�ŏ��&.{ܷZ]��QWt4��l#�K3�Uux�QKF�xh���)E�H��mcrj�{*��B��}����k�6WQ�9�������
 0Ju1)#>k[�K/mF��i�`�����=����c�{�9׆̓72X�Mr����[v���AQ��,�#	f���j������*1�ܘ���9�{Ӕh���oɺ�dX��T������e$Wf!�Z;��
��f�+Q��N	!=�w;o�(=�H;�6\��mi2��T�J�Yq܏���C:(Fܽ�-���\1�0�js����d��7�u��̬W�4u�v9��\�(�}�*��>#�`���Zn�p:�D�|�	��bH㞼�Gp�VRԀ`ZI?�Ա�)�U�~��������w�
��9��=��Ջ��A�O�w]Q��/�̙z���8�?,̊#+?�������O��-���Z����]+'H�q�Iu�s�j���P!��^���/τ�ެr|�#L5��'B�"�4��jɿZ2@|mpD��|�p�Eunk�^�%
<�k:�(��l	n�O�'���vr>"�HB��c���#��[�2Y�ߚf�GC˦�� ��6~ʂ���=1��(AW¯�T�.����Yp�k�>�l�If��-��3��m-��ʕs�B�� �)�ʞ�F�68}.%d���/�h��NM�@�	@��]RLSUAH�U-�شe��Аm�qЪ&��c��1�%�G��*����qwhP���z���:�kHu��4h��Lѝ�]j��)�i��ۍL\A2�P��	뇾[v�8�Z�z��"ӆ�U��=�Tg0�A
5Z),Aߩ�aDbI��,���⃭V��B}p�l���L$���m��qL���x�X����槖!ٛO+v���?��Υ��_te��B�x���?�ƋdK��N��]������	��uF�=1.^]���?}u�����d�l