XlxV64EB    fa00    2df0�ֶ��H�L������X�a��E�菃�=%�"m{��8"���.�F�Ua+z�x��Z��7�4��#�t%.��n>r?#�/ ���m�J�4b���Q	r��o�"Ǹ+x�`!����B=R?R=#Q�A�+}�?�	����	������%����o���(���⸦���qj�wI��{UX�:���~6�&0|��Y��/=7:pT�W��f{ȯ��%х[���˒y{yR�楾��2(�w�_��X4R�d�0ݷ>c/n�t���Z�_ȼ< O��l#%��4z����uYӟ�\�&/����V?��tM���o�I�+@/Ֆ�s��a[���[Ԉ2��`]��� }��$��}T���	��E�L����?b�%�a���^hl�����/�>�U�@`�����ea��?F/gNU޻��ӈl	[�o[�`2�u0�ܴ��B�gy�^��	z����
'�h�J�{����F �u�g\�p%X����!x�E4��cۏo:Jl�9�%(8&U�Kj��9��UbS�i���q��Q�����[���u�E��V��7�:����2X�6|�������if��T(�&Ѩ�f�.Y��TH?���
l��<�?{�w�f�A�����_5[�CV�\�qȊP.��6W�Ⱌ
�96�W4�7�'��2n�V+��DKs�u��7�������fS|Ï'j^��]��9�W�*��?�/���5"J��-���K��5��5^�����+���G�ȱw�p}5���^VVϴ0�h��?����9����ҷ��f??K��^�7Ê�];<�f�}*��[��	�����
����W��﬽�<cP̏��
�S��p:jK^�������RUL<gR�r�I�[% �H�a|�����Y�C����%�<h��	�!�W}��4�]d7}���4�@P]I�ow�u	������s�!\�����V��,*�U�Dz��"�K��椟\�2�g���{2����x�O%k��a�Ye�}�Uoa��t8�&F�O� =t��[��ޚZ� ���	�r���<�?޲a��V�(�]���'o�Y��@M�� ��t��02ƚx��	�`,�7�i�#z�F�ë.��J|�}�`��:������c�)z�
�)���#xa�Ar��K;=_�r�r��/�\O����R S-	�R՟��/>�| �:L��y�����a��XÌA'�Iu��o=�����ۑ���^����sДQ?r���iyð�f�̘4�<Μ�7���_m�З�	�D��:��CEͪsWq=C�Dx/.�����`L�����¢��>}���5l��H���^�VP�Y�uv\g��,K��3:,z���?su��r:{}l@0ߔؽc~��u��~Q�<��eV	����m����`d��I.(*0�4?8x,z����-&��תcǞ4wɽ#����y�:�]�5�~j�D*N�&�O�>�n�q�j;�=pd�J�V�#cT5�T٥E�KJ�(a[r�|Pyūɻ�$�8���Yq��<i_5E���Wɱ<Ny�j�oc��y4���["����!9��	�F�7�ǯ�׍܋6�u����5�!���J��9������d��v�i��:����� �J7'ް�\ӻ#��5���Y�J,zp�:��t��p%կ#�"��_Pe�Y����-��^��m�����'Mh��g�$hG���Ӧo��Xvo^�uy��	������<�n�MhU���s1�s�Gޟ����͐���#a�)ݻ�P6��
�KK�E��Nc{�����>�ˬ��ϼ
{Z�}�s�Ĺ���&H� jAͳSA�Y�d �J<�F�~3�u�+�+F�W�kx���~+Ii̷i)��	`7̂�[?�
	�&w�R�[L��21�sC��'f>��־?���č߇?X���$:�?f��rU؉�~М\�Q���#LO�2PR �b��(���Fٹ"Rm,~?y�3�����s���p��g�^*! ���A�:E�D:he�!,�#�1�,e�:.�h�w�Zc:�% ��T��y�S@�}���h�"^8�x�[�~�9�R	e��r����@_��Y.�f�65l�*�삢���#�����,�?����`����ַ��k�� ���leC�u�+��i�I�Ҵ�<ٝ�!U��5�S|Ԝ�f���g��m���1�a��Z�¬�5��3`�82>u���g���sJ��<̣�Y�S۶W �.7����sN��T[7��-zn��{�kڎ�'h���W�W�;Z���?�VN+��'Ρ3X����l6�[�G�;Et1X(V2���y;���7���Zd�`�� qGX�f��.X�x��@-cEQzG Sk������w=G��q�b����
��Rw�ӝ�ڻ�II  A;2��İ��%VM�3��`�C��9�\�d?�IΙq�'V-8�t���&���dL���[(	%]��g�Z����  �2�U��E���ea/��Bc@�����>����	50cS|Ï�l�~ɠ���/�h|*���T�ה�G���5Wr���>�Ԏj(i8h����u|%�������z%Ϩ��qK�� K-�՚�����EG���~�Z�M@���e)�N}}}��$j1������?p"x���Z�*wӄ�Tt�&۞m��f����QЄ������ЅS�L�?Y"'��ޚ�¡{&��#��sr�(g�mG��!��9|�y����F�����;t]m{��m��I.jݼ������a��[�H"v�tT��ҡ���������ґO�+��J��1<��v:K�gz3�h�<�/,��"V𦭧�޾��7��a��E��j6�Y�9��UM���\���RxV����&��}��XC[/CS�L�a���2��LW`td����b�\#���|b�T��n<�5%�e�V���g(�u�r�4-�E��-B���0_]Yj�ݱ�d<��b��\6�??�x_,�a�?hEj��\�8�a��C�̉���{�5z<[�Xc���ǥ�=ͦ�x�����d�:c�X1��td��c�!e�B34�`��1�Q�a/;�}�h���si�]p{��������Y��6k}P<�mpg�+��1��`qV~�[˨	y01�w�0I56��D^�Nu�`���W����+�zݏ3��ٵ"Gr�zlw�ZIq-w �(刀�XI���g�V)���T��";���w��FB��9���er^i�������ߒ�Xh��$N^�b�
�L3��ϏA\d�dQ~�p2H�E8���*q���$X
�6jyj	�_Q����c�
K� ��5�M	�t�
D������)���l�s������Ft����l�ƦF)�0���QĒ�a�ڴM�1�S#A�����[dd(f��t�����b[��0�w�W}K�+z�du_�P+�y��髧<����j�.��5N��mpZ�M�MC�����/|K����.G'.F4��󫳕έ�����<�n�"d�#�B�6V�i
k��i�����+d �p&+���]s�$U�T�[t��k&qM��byz�"�&]q���ÓBkS�^�S��Z�fwE1z�59u�����i]��ʞU�M��:v@3�`!
��4�)�,\��$���K�W��w��zDڜ;$�L:�'ԎDG�ɗ1��|���@����lW������@�\6�Z��}Q#'�����S���;J������7��P��C!@\A�Ho6Ddz���Ʊ�s��KU���IB��	7�)�f�l�7�\��w��9LT^_���<���5�SW z�ND��9�1��?��Q;���O���@@����ض��C�q��SB/����'�?c�4��z����/��jU�����S?���Wp�b�;��=�r�	95�EPm��Rȥ,�j�:��8� 2ٲj��F�>�@7���<��8]����'�9K���r�%/������v+;���0��8���e��ze�y���0UHm���;�vo 9h��O�
�";E�[R<�M6aW9aղ�'Yv�����/���(��6��>������2��B4?�7�P�����(�����Fb<�a2�#�	�@�m�4[z��&!��#���oQA��/7t��X�Bd5"N���Ekq�7J(+���L�7�����۪9|���W,7�f��r���\{��L1�,�� ���!7��U�쟱K�G}����29��ɛ�r��{�V躴k�"G�]o���q� +��>�4�a�C+�v~.9�ʟ�lvg���ؒh�[�1�������ď`j]�|�Mr��ܿ�v6�]ϼ�r�� �%b;�B7f�6�PB���Zi;��q���T�w��/���x��>2�4D�6-Ĳz����a��h���|�+�w9�$� c�!��^�5T�`���>
����>�}�L�Y�Y�G��Yǽe���&�6�Kp��7� �B\�EF�#m����)f�_�z�nt\3b�Q�ji�W&�6�r���64��_!4���N��p�O�-���hqE3�ڭ����fc��r�#Ap7@~IM����h"��<��7,�c$���������Y�8���&���2@������f��g��̓}����نu��CE�ӆj�$u���ZQ��3����c���X�XO%?�GƮ�ם
�D(�5���=����~�:�����V�X �q��
�����N�4��ZY��عF�\w��]�F+���(���CA��5᠐>�	P��)�����΍�q��:>\802����8r*7��8�װX(��;���7Y��d9���4v��W��b`l��w�x����M)V�n�j�c�+����8���0U_y���ά}H(QH�����K�@Њ�k�XQ�e{��xN��GS�� ���7�I#c�Xʈ0���P������������R�j�I5��MJǴd����4 s�����i�Aύ�Y���N�L��hy6c�Y�xc!q�hN*�(�GEX^����TʔB�xA�OlـDe�)�Jp=h�w�ےd��5W]�wx��I]�����js0�����gyf����5Г��3�	��,�G[9�3r�3���oILi���yR6�亴&�������R��c�wK��i�|�ci���"~��Q~�.�
V�GU�D4����wW���Y4nq��"�^�Ȓ��%^�L�v�����r.�����O�Z51�׸������&��D�=-z�uu�<�n�Jz�v�cp�u��%��+�JN�9Ùwf�qRс���b7/����]���7�@��a�#��Q^>�<��h�2��-8�@Һp�(��9&l��`���C�<�Me>v�mR��K�A`��ϋ�@�^OUݗ�#��~��|wˎ_���|׽�{o#�{���� 7��S����#��%�@�ᔧ�}nQZ�Q�'�G	ɕ۪��M�����&ߖk_����N*C�t+"�?\*d̵q.��$Q�5�fF����3m�.]�=�
@���ኢ��#Ja��Z;�x�k̙inAO��Xt���k��_��Wĕ\�* \�����V����_z2�X�Fq���˶�)���/a��%�Oܮ�;Ft_.]�ʦ�ҜE�ۙ�u����Y�I�7,'���O�a�/�n@�i��,�Th�x�U�����_o��Q��h��b�ڑGQ	�*�����j��hݭD߿�?&���*���i\�g
�U�#�� �2!�EvaA���)'��:�9��e�BB��6Մ��AL���cn�X���bN@���]r0l�g�X�����@��a7�b-�=Ӥ��k�Bt&���]����{��U�w�N҂��=	�q�ٮ��`F�z��6t�`	����`�����9`�\���8{oGQ��q�1J�}�~}K/�l�ۼ���9���ac��#�@c���hէW�i��O��dmof��/)o�Xe4UU��{��W7��3����$P���Pf�ׂHބ��ɴ@L�%g�32��߹�D삾	��^�M��""Ķ�b�qVZ�iG� �&����p��K;��������Ѓ����=�=�oID���*���SY�E�+�����y��Â�#͎���9�K�<��	V��2�zV��:�ȧ�5��]6����
�Qsl&S���,�M��-b������R!��<��|ceA�M�ÿ�\�갸��QY1�{��H!��]�^u��WJ8�$�h��@�!��"(�i�C������d�B�1��-��H����8�xM�'L��oǉ�<*&h5[�AO�Ԃġ��/C��&A�_y�?�����lq��>GP�^��k��~�p��VE�Y'�][|n'A���})�닫�d�����x��CDag�
L7�3�Vn�ݟl���k��)��il)5;ے7�V�J%�oH3�܃�<@�}��5�}��Q��4�8��(��>_�
33�c)�8��
���#,���~LK	SZ�Z�1	�rm�q��f��Ч�jA,����̫q�!�w���,���������jQt�5CE�Oà_�F�l�N�.nYtv���t�}!&�e��g�8$u�삸�G0=Mmk�z�`���a8�hn��^-4I-t��4��έR�	-�SX
��J#���B�T��0���EA654)u7�j���^U�?�#l����כ �S�������[���_�7I��E-6W+�6���w�=��=W��	2z����<����R=;;�@�����c��."]�>M�&�3��D�����0�k��Y�bǔ!hD3�/3)�+��'�����2,��t�|߰������%�̯�?��� H ��ӴO���,��p_�2yA������hIm��|��][W�+��bZ]ӡ	v���>R�)�>�)p�I��i�+�
�%F3�	�pE��l}�:~1�u�������Io��*��{��T�M���M	�����n��H�&�-����U�D���U%�ʷ��
��{8��v*P���ؔ�9ֆP�1�����g��eE�˜�{M��.�Њ%�]�u�'=��� \ޟPF�Ȼ�t�ӳ�k�+�oo�H*8J�/L���B�X ��*r�{��ͻm��+�i����4�NyP�[�!�n����Vо�e��������-���	e����9ndDXty�� ����[�=��R?>X$ͫ�KȽG��X������<\���z�rO��k�;�~�Ǡ�y5���w�l�0�s�G�\�Ǽ����d�h���2�,�RB��3�Z9���"2��A��)u���gZ� Տ�*�F���Ё��c�o�7*k#�P��ͼG�w��z?�a��\��td�Bs�g�G �x�~�HQ�`���Ր�����E���b�gU\����_w��A�*�������-d�s�Ƌ�2ݺ+_��cCE�&�Ɏ�5�ϪH�x�/�jp�R����4��j�=Y|�X��7�`��
�d60���"t��_lP>f>�"��a��C\"����N
٩�
)���;�w���������$P�Y�́Ɔ[�3�!�p����bgI[��1���O3��%���˻,�=n���dB�n��#A��G"��S��(4���9H��ޣq�Mx�ұx�(�!����dVp4��H��C�B�ܮr���}r%`�
�ƽ�2/���&cx�_Z�΄r���v��)D�W.��D�b nߕg8�0� ���5������QJ��?@�M����~;fjD���ۦ����Bzy� Ì�����hX�����t��U	ҽ�W	�H� ����e���`I��1��.�'�C^=E�KxAT�G��=���ψ}d�t�DGJ���r/��m&�]ꗖ]T��~�V�W{�C�i�YIQvW^���1�B!"49�2��=h�/&�
"�r̫����+�VV���1��!����V��ي��<�!a{+�[���rq�y��\���^!��^	���u�Eߓ�m�O���Lc~4�}R]G�E�a�M������@�i���^�¨������0�)�s����\K�WH�Z�4h�C����c���z�×ب N�(2$H���1��՟��gv���,�h�lN[U(��ƾ�
)����N���3����q����x�([Yj��Z"X�*��u:��x�8�lo"f�hn�/v��q_���"�̻DDv�����.�C� �����QQ�w���(�jǟ^9�\əJa	��}_b[��-��G1.sc��ƫ���Vh8�S[յ�"�E���/�3qϮV5޿�	T(B�d�x?��z�H��?�b�j��������rW��E1�Wq�ZC�,��^W���ﰒ��U4��!^ @F����cL����ݍ�V?��I%A�s��}��k�F�`�+�U�&�g�7y�9�����
��'��%	�Ak%����O6_\�sSZ��8��*�Y��E�.�cDW��"?=�)�Ņ|�G�,B?�^K�4�1M��i@T�2�B�f��Mi��F��f�Ņ�5X�R�a������l��j>�

J�N���	�vZ�ə-��W���S.�=�m�w��9)���ԍ�h�F@��ਿ� I�B��@�c��g/-fz��O#R�\!��]?D�P��-��f�l�miި�+�o�vw\׵�eZzmL�H ���]ǧ�}����PضoK���	)9�B\��\�c��6��X����b���� ���t��´���7T>�߼E�S�
%�g��${�9�'o�[;���Ec� �jJՃV�&�b�"10��-���5�Q��Z�GG`g[N��癥o$^{)�xMgal/q���z4s�pcz����w��Ica���ҿd��m�	�d�C��{���0���5�L�����$��N��J�Y",B�w�}��`ת#�J�H��$8���I���o��|7�����������8���w��X?{�vP�cs�����)�y�n)��گ/�Q�9�p5_���R����XX��`8���٥D������s�gv����ٟ̖@�|6�־;����	���W���)�i�\P�Rf����(��Bo��y����î�Դ��e��[�n2٥a2�>JhJ$���=����Y�=5F~��P|��KP���r!v�Q��餇��h�����5����A�s��$lk5~	~C'I-y�@�.��*K�
e��WA���m���c��-�b�JÇyŅ�����p7��C\��mw�d�HAER����~L���7R�W�*tQ���,_$Λ>����ՠ�`e��&Ck��yHŖ=nle(����z���	�J�`�B��z�SI���a�ˡ�@�w�Z[_�Nu�k�A����jT��Y�3��ΞKcYz?��A��Kj���z�FE����)0ْ�r�c
����=�)p�\l\�dW�����;Wa`0�iCS��و�t�Y��x+-E�{f�aS=4�}j��4�\9����,ˏ����.�yE����V?����a�
�$�-���gz���Z��4��2�.2}iE��%�UBE�7we6�9t�E-�	�m~d;����&EKʄ������#��{"����d��t�l��9W<D�z��kQB�>��\73/k:��	�c?�n}��P�h��gK�x��@ܛW�%3p��#wε��Kd�)�c�&����`�5L�}�\��+����[ ���ʲ�a�7B����XZ�J�4����\��&a�[!�c�O.�=��洔�Aue%�wV`IМȳ�Bplޠ��]�JS�R�=�+���_v�x;��/{i�9�#Js9�1_r�4P� �V?���1���9p��%0�[
�\�9Q{�����kׅ����㩦�܃Zf?3�:h�
cɰ)�8 ��	y-�J�r��A���`��$1l�a&B�U�r�e�v@�� [M�cSAS�� ���}�7���/������߇P5;њ1�� ��[#���x�40T�7��\��Yky�Y��6��詁�NKϫIY�Ԇ{�)}6T�ҥ��Z����ߥV��������_�I''®�R-F��"���+�{�;����V�͘y����PR��S� 8��C�	s��OJ�[�@�쫽�ʹ�(��&��[y��n��|//.��s�v�$z���غ*�/�n5�7}!�=kX(�g\�����fe��ut��x�c�t֝�Fs�i*�:���[Y�Z�5;^J�����W���(IF��0�=�-l��W�Jǐh�>���?�DK{Cd]��L�m��/t�8�B]�м�v����
�Wh\
�h-m����E������l�gf�|5�!�SY}��΅�E� S����crC)Ē�(IŚo��x5���Tt�"�#wJ��n�h��x�}f[�~rl �y��P%�uW2���"�e������
�5���A��@�xv�) k��<8[�1�'���t �р��j���ޅG�����{~��+7Ok
g����ɸ	��DDX�Hl�&�n/y�K�Y�11l,�!f��\���v��ȥ.�Q>�o�^O-2y.�*�0�]��x��c�~֧@.(R�!n�'%1��;�_Ը�u)��O���6��V5��[v��3:�U���*��>�=�����'>�e�d?�O�a-��߹�42�)S1>��~92�:@���-�R����^�09���v�n(}l'@�(��ܷ�k����E�
3��2�2q�un�2�� ���Z�{;��n���w+�/��ss��/�Pl2��[�}A��Z�U�$�=���@��T#�d�(�o�>8�0��C�Ѓ ��%��ɕb˺��1`��" B`;�:>ѩ��z��M��W��aR����/�6ٮ���
�n��?3��Q�l���-7��o�~SB{lE_�u�8��L��Hwћ Ao��S�t��o��zw���}�ct���giY�*�����������"���+{o�3cz������{�4�+�*�*���Z��P���\�Y�C�I0$�w�@%p��"!Y��aT�Ew�#WX*��m�����#$g�͔�y3MP��l�@N+#Sr0`��z��{�M��Y�l�1�F�5�����h!�p���,�K�fq�ܜ�Z{
�E����� �/� �y �le������aTa�R�Q�#]k�x��ߣ�Ę���t�$��x�$}�J8C�Nb�`�s}��;b\��â��-A������t�>�{�>��v{#0��nxAӰ��z�~F�>���Brc�B�X@U\��e��I>�M�d���K��!rS(��>o���fc�ʗfꕃ��ᡣ���0���e=��l��k��j�vI�����6�U���tl�ߺ��pm��9哓�8> ���lN��[�)7��A�?�o�u�U��G�!��Rz��4�[�G�A�v�IE7-��V���\��ht^����{�[������-�3=�;p�`��� �⛑}ʃXlxV64EB    b349    1b50w�\�3�i�섴�r(?�h�%|���۫hA&ǻ���q*���E�p�q���f�1�.�Hx�vF��+����&
3��a���.�U(��M�<cm��VY˟`�W�$�`e�����' 2����Q��.��3ߐ
G���[�l/'*t]�N"�1�&��{Ui��x�	c�3�-�M�ڥ���&�W�!�A���\�5�7f�I�f�����˨\Dhۍ�%l�8_���Xŋ����N;D�gaZ�=m���}޴��;}��b��mJx
��%�S�l��Ox6a��1�����e�y���7eo-��#�s�"n�)yS�GS��S�lctQ���D�f�����^�]��>�����ŵ���Mq'����K�1k��DI�ԧ[�Vďa�Rm��*�O��Sߚ�}�<1�{?��gP��7��e�GVT��'��;�kj^���U�#�u�1�}(��$Z��'���l!Y����@�TKL�tHC�7�_P4�I�i��|p�d@��g@���׉i���9�����Q�A�� K������J�t�Cos)>�&��r�.���M��G���Cn�N��9�o)UQ"c�>����S���ܲ��T� ��/��	���qC��?��`h�cj��Z毓��QXL��������=Q'������Ͱ�#RR`|��f�j=�,%,�Yc>P `����wB!*\����i�O!��~B�ɀ��I,�eK�V���
�w���7c�e;���c�/���'�26���֑�E>���>�� �E:���Pe( |�o�h��:���_PSW�yץ�v�6�skt������r�Sp��w}�!߮�>t!��4}�?p���(s�k#*r'����_[�ISEn�&#���T��L�@7ކ=����I�b��'�_Is�+�2�m��'�9������5�5m�i&�+�#+s
�*��6��ƅDJ2v�y%F�ƭ����������-kRH(�%�Dq\��.Y��e�/�U�i�����^Ɛ%1��(��H��^��ۺZ��O��)l�Z��X�cVo]�l"z5Z�G���Q��&x��~Foq�a�"�ps�(��PbU'L�Q���3]g�����z+�agD6i���,vI����!ߨĢ�d�s�f����>�t[(6�>�J�$!kF����&jD��zbh_��;�8{?Dr�Z�Tz�ye�O��~�3�T�y��۶��R��>��{��{�L�˻��]H�y;]��瑶�J�,����a}�: O���f������ӈ�5Q��>���W�D"�Dx�zR�H�>�=b(#nER���H9BV1LU�LI21v���~2Y]-�@<0)
g��Mbg��?����T�����s�b���J{������"��td�o���6��hs��WaS���;2 �ꄯ(�V2���EJ"t����h"=���7W1*m��?#��@�<Ãr��>�sl3�L����`�U���z yms2����������6^>Yin%~C��lD!��=��TGo���ǃ��[�D�L@H�&6w��G�M�H�x[�C��P�����	���`S��`g����T�10d�����J4�e�����]- �4��� �gJ�o�2ġ_z)��C5J�π���j8Q\��h���m&ߛd7��;�@�*�bp?b��9|�ҧ�U����iH�
p��|��Ɩa�N�=���'�{Q�Oj|�~gY>b�?`i�����}�:�|�ջO_O�5�w&C���O
Ć�z��|v~	{�#N�
�`���%q�����Il�r�r$8/���HN���~���o>���Vh�\�(J7a����V��q�U;��"R8���P���/�^-���ޒ�������&y�Vt��R�^��N�y�( ����F" ���"kJ�:�]V�¦I��1��j�F�HKL�T���aX�1m������ވ�e����\�X��G'�K�3�|��I lE�0�\*5����D]C�h�=��M�Z��G�K��)W��+����i�!���ש(ŕ���>u�p���24 c�����
��騑%�~�T�/y΍�Ȝ4z�;���Ԁ�G�bu,�%���i3�ª�
A����iq��1���@2��;����j�Bxb�2�����;�`�r�������rS����u�gqX�9���8��-jE;s�d�Bѥt�c�d���~"�x�
u#���3f���c��5n��-#���ݐ��G(v�-���#��!�@�k#�'X켾W�'���:��<o��8�Ơ<u��ٕ1�����n�TQ5���� �����3yC�xo8�W�D�(p}�&T�g�GtF�C~�YC�R�`T ���6��k�~rkR�d@�cu����j�������A���W��� ��ܸǦ��Dx��G�^W�n�'���a�u�����N��C�b�=�l⥤�L�Փ�x��G���W+�����"Bo��*;�9u�SG��PZ�^�N���b,w��'J�:^�2��r���M=<�޻�j�U���VB�Ji9��7�A���PF�'�Jx=�T6�@f٫�E�x�A��ɁT^x9�Q��j7������S��O���ZPR�4iY�}��y�{<c+�M	�k��D��^�q������y6ϞRm6�<��<�	d#V3)��dF.�Z�͞�y$_;O�/�*�|Pq�N�,�6�?���G'߱�lq�A6��D���djO}A&.·��1p�ey����~eL��y٨�S�wt@1~e��n�W	61�Pb�[��ݺ�m��7�m���J�	-�X�<Ug��z,���*������>�)M���+9�t�b�h��j���m�c�%o�p�jbI*��"�$������ �_+x[�w��,[��vH��h�:�z����z,�Uɜ�@��%+$��#@�Oɏ�,�l�5և�a�'�-V��RU�ݛ�8t�(�+�YN�/��+�U-�nD	����~'PL9I7�=������sԙ��
l�0.�/��� �e�#T��Y��7�cTLa�a�=�Eo�.�W�B�1�X`�dc;�Y��Eۚ�(9��09��98ґ�	:2-b��
c6�l�	Vs�^u�%n�:{k�y��&�z����D�:�Zaa9�e�A�¼ɣ �3t�\
��A������"���Cy�ӿP~��Z�]V��	4O?	��vn��H� ED"�ܽ�)�8�V���?p*���|����N"���a�ޫk\�i_̞_���8�v��t�o�[7�g�`���09Y��nB9���Y�B���Cg��������ץc1��q���E�6>��VU҃�;r�!D�H)"_�3���9!���o͒εט����$OzȚD� 6���W7�mPG<Rnή��酎F�,a	?ñ&EqH�c�T��S�����h}��+;���8��:6R����(D:T�2��m��1
8Y�c�f,�ǯ�X�zF!T6#����v*�Q�A����i�[�}�<��>��R�sƤ���*]ۗ�f��{��K�d㫖�x�|�YXX&c>OF	q9���:8Lj����q~f#nf;S-�@S�4�PUd5�%��DZ����C���B�+�n\G�4 �9�G�	ê�Hʉݍc�MqىtpA�����`"Kt���g�Fԥ�rS��$�AY)�ă��S	uEIo� ��,YA^��[�No�~6�U֠�AJ��Z�~�+��q���Bp��>5����{�حk��jF	Ӳ~�4��'e��>���P�5ץy��t�@�ڶ�N�&�D5/����W����g�>��𚀗f�
�����l�a�t���>Nq&��!ŐL�?�PgJą,��&���P�kh��rǫ��*N��_u���@P�XlY�3���j"�XM��b{���I蛭L�㐌�ݰ�7�K\֒	���m\
e�{lqt!��4�/�[���oƯ�T0~�U�#͵����uc���Ug�trʅ��?j�X�v��z�V=}9�:nݺ�7�'[�	��[QQ�>�`N��j�Kй,�:R�auJg��I�r�'�W�؁��u�)�����0�i����nw���0�y��@� LGմ}��F=-#�y�(��O f#�K1՛�|�iGt�����|f~�n��R�UN�=�*�W�x�g��t!&Smh��3�,�L椆]�!S>��?"�.R�H���7P�-��J�չ��~����D��Q����r��y���ԍ͟s#U��`,�.��T���7ψ��_)iߠ�hD�-h��]~tG�n��T��[1����\	�F2ǃ}���1�KE\a����IOخ���V��Up^��)>,�$;
�I���g��.�V>o�Ţ+f,����ٰ%����9�R�}����G6�U�������ɮ�q4��!$֡xb�)U�Pl�?`k��J/�X��Eh�vK�Sn���;�"'P��'���J���:(~�V93"EWBNN�X*��d���2뛙j�d��i��;���x���$�"Y��qu!d�+�x�kj���Q/De#�Ǡz-b�����t��p|��0C�m��Fr^�Vl�Mg���X�Xz ��;��{��S�Ψ���%�5\:)�N�4ⶅ짦�������Z���Y�%dk����s�T��d�}5�3-xd;�т�B����Mʚ��KI���`��\�ӣX��~�����9�+  )g����uM3t�Cāq�Y�$��):���O����]��>[E�)y�;�:_V�)��`�$�A?��H_�����DC�^�E"��4�$G� .���/����Nِt����b�H@��G�x�y��o���^�ס*��R2�C�k�_�<�G��h�Z��,0V����N�ʅ�?����]|u�����4�E}�먼V����ס�>A�N�E����_Б\r�c��Z���.�������vu�ֿ�	��>+Z�*��-��.E��5�����/v,Bi_����!������^�7h{2���nF�-�
9� ���6|��"}FغT[�^8�� �}��98�(�'��%̝&��sAQl �E�v+,�ܮ��1A��o&W��`A)p&�|J�Ë��=u��h-�d�>z${_�i̘"K��AE�j#a=������(�Zwؗ����%�K�zX\[�$�X|�
M�����8����x`����獄P���lMv������azGS�Ir��̳V��R�r��{�|�-�b��������敁�Y|濎��:��3 b�8�w��J)��H�w�;�8�bj�o���Bw�P�hgz8 �l!K��-�@4�W�-�+O`o���1d�t|�T���<Y��m&�1�x{�5����9V�J}-�_C���]�<���b]���^�t�X>D�,�A��.,�k�D�><!d���E�c�Y�4�������kBH�F�ġ���J�v�1�؀g
y�=��ɻ?��d �E�v��xc��"JN�U�X��<��ŒWq(��S����W;�!�	]��7�hZ q��WA|���}�76)C#+�w�|r������JT��+�]s�bۑ��_�u@*{���Ӹ����-��$�.z�P�yQ��0���)Ţ�Π�fx�N+B˙<b�ga`U������9ja0kJ������x�N�V�����S��溦�WCi��+w�cw�&�~O$O���y�����J�XJ�GӃJbR�����#�}�ЪC�뗵�-��KW1���T�*"j����ɔ[�j�z�^��"�Ш�'�o���<^�t�$�"�0�����'f�G�.���p�##|2a���w�s�ÿ�1��b,�G/bʁ�P�Z��Z�Q��.ok�I}�1�:\Z#s��ދ�Il���g�\2��3@�N	��e�� �cb£YP|B~������5b��_d��c+R�p�7^O��"�?%q�X��K*½���=��� �g��VO�<�R��1��� ��?�x(V����a�?*U����e����hh�X�ob�n\ˏ$[O���/�mW ?%Tb�狶/At���=N�C*2��|��ZZaޛ�%h�3��#�v8e����j(.�J�rJ�ܛ��)��6ԩj1<�Q�I�Z����h�x�$�1<�c[KKA��^�*�?
�iw;�O�@��Ɏ+�c����9���U{���_�E�ds����F3��֠��X���ó�Y���af�?O��O>�k_B���P�G��|�! ���� 01��\zG�XzF������T�o�'�p��6$�D#s>��&f�[�G�t�+��� ��^a�j��(�r{���7d
�r�f5H���Ҩ�&��/	�)x�<�I���=~5 %��+��ٗ�B�6@�b>P�++L�o6�&�K�͋(���ҌEa�@_2KI����5^����6�f"Qm�Fs��Z��#��Eˏ��y�2��Д����H��V�Z`��J�2E�{,T�Y9B�J��ڛ��S\���V�t$�̄kJ�Kx�w\2}'}G����һ�l����<A21��66)� Z� >6��ye.t�z:.5�#�,����%����>�IW��y���܇�#���GJ�q̕28�;QӱTHJa�`:3����a�l�[6>ˠ����`F$>�Z�Wt�_�����4fڈ�"�mwq���M3��,v-p�_��������c~�e�0�./����5�\��`�	^�	�ڑF���?p!�"u6��hXʳ`��;���7���@�`}Z;'D(t��4d:��(<����O�
��������"h)��$0�