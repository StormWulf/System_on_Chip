XlxV64EB    182e     880 ���ƨB�M�4�v��Y5RL充A�D�7�4�xW)�MA�{�H͍�����6��Ԫn@�;?�\O��U����=s�
�8�E�s�(�<F�s�]M+��"��b�}�G(b�(ϡc�L��>�������/0G6�D���8��x��.3�'���q'l���!�J s�s�>0k�U��Yg+f$�W)ܲ�o}J�f	HQ�|�<?#��텺'�i������8cFy�'��-�˗�o��޼4����w"sB_��`���f�����'�+T(k���S�.gf;M�h��OA�e�#���e�QNРo~x;��Z�}�� ����Qb�IV�M���Ÿ�w��v�%��@\	ˍ���D�.ov0A ����p?�_���7:�0J��uɓ��|os'��� ���wr`Lq^Sխ��h���^8����/����@d�[�6l�P�p�u���,�;�h2���#r�H��s��6'@�[���*��۫�v�`㧄���^ �܎�k"J�)h��K�vP�f�km��}��~[��zB�ӧ��|�4��k3!'4H�Fzyĝ����`]=�O*��z�z�F��lB?��RgHƢ.�I�$��#Ro�X{��Zҕ���2�w	`5�Ydi��R��l���X��g��Eb����Q�:�P��������ε��О,%}��XvF��k0-�D����KZ���9���J��"X`G9��!9e{��F��0��0���Ӂު��;ʌ��4�����i�|MC��~�w��@�O!Z�(��ϯWa���Lro4�n���ͷ��F��ZJ>hu��;�/���>;�9r�a��ݧ�]Ё��LԺz�`&��j~��y�X~s��H����_(�a�vB5���թNs�1�Zn�B����uA4M�4E�� B���̧������~�C
*�� 7��@%;���)Ղ�g\gc�K ��-��"�鏂���])�����0@��`u�\'A���:��T%�f���pNj��kjD�R�A1���I�΅ˀ��S���CO	�^.N�����X��.ظ���90�r�������A(2^��i�B��+Ib3+�,z�������E4r_�	������T�i��H�N��ҁ�f�b�f��|���FR�Y*�����&��8φ%�<&��@B�*kt%�6sF&R��.xW2DO�����Kd�Mٸ��iQH����3�m~n��?����)��;k�!����_�
�qr��}�]-uc�� ���Ta�gk��/,+�����\+Η�]��d��´O+!�-�vd䑦l5v�� '��A�B�-ٽ��L���ųj�و�n�YZ�ݦ�U%�,��Q��~	�R&��%��gIڦs�\�+�¼=Қh$T1�)�Y	m/���^�`{����)S o¯3�����K`}�%��>�Y�i�&W. "�zf��╎cg�RT�g�0vv������ٜȸ�]�%�ܠN�������Ǭ�����y��Y�Y�-rO��x�[~ř{���V�E E��+�9��W�������Fqm�����{Y�2ecaШ:C.��Wێ�*j_K�
[I��v�!	)Eʥ@�{�i�g�ã:��Pw���D�U�F  �3� GO·#�e}�:��C$O0�U!ZkcR Н*i4��k�F�|�k�O��%ܤ��`b��.J^��!��v��`�9i�~4���)�
, �	��>�MN3�P1��T4�7�$�*����1�i����&0���xN���ڜ��lE[0���`��	͇�wi� ��9�-�ɂ��0�"戯1����`g/r�%W�b�m{+��q��:��x��e>���U�#�sZ��G
���F���d�N��q Qm`hҺ�35�\��i�i����{��}x���"#���|_��=cy�2��ȱ�MRA��r��X��O��	��Zk��a-JaH3�L�e�9t��Yޛs�� ���w�y[��ځL{s��-Hxb����
?�r�(K+fe�5�0ps���2���t �32���߇O�K��W�/�Z�94K�d��5q���|̉b9<j�!�FΑ'�l�"����T�Αng��~:O��Ⓧ5us�