XlxV64EB    1fd3     ae0�,Nƅŗ^�I�̙�I�'�y_�&>�%w'a���$^|�G��a����{��L�x�%�]}��/��Ϡ��hH���2_�A/U�#�����ڞ��`�#��R�ա$�i,�`�zdXs���,��@�Ү���%,���1�%`���Ow�����޳5⋒O�<o��~�U�G�\T�l��=Y��F�I�L�.�*}����=L�tI��f�a�'��ގskgʏlv���L�Y��@��<������}����`�3#��:k5b�.I1,���� T��7dT�	��T#�>⺖«	�o��wn�w-�!ǋE�}f�@�u�y�BK�����;��'̈����ew[?Ɯ��}vÿ�u\P�f�
Wt��tWtx0)��pT�����.a�0G/�I�6��`y�5��:(,)ly��-~��7�8�*t �e���m��V/��Y6�%.8k; �q�/|��ɳ3,��4[ȦK��@��N���3����g�~�
ƴG��a�*���x�v�?;��|F4�����G�Bg<�	>UA��t� �Z�;�I��2����k�='�������@d������Li�;�k~��x��O�*$:���I��UݗH\V�Ѭ��?w�.��q�l��u*�iH,�x��dg�4˾��@E�_�=SW�H�,���^J�XU�lk���u�R�?�m�o�3Yv �Ud,{ �o0�Bo0G8k�<���+����C����d
dU_�i��j�n%l��y�_����@��4/��B�w���5$H���m�+�أLj9^�}���Ny�?I���I�~�͡�^�d�t��.Q߻1#Z� ay�Qb<�t�A�bRc���x��{�b/0�?�g*�#S"2H����玗�Fu���Z�b���b.�|���Iu������2�1��'@y{�KN��|�o:3�j+�{)O6XU���x�ܰR��=���&u_/�֓��8;f�%( ����L����uy���.WhLR.��a��@�.Q��Q$�����V�f)P�.[R�xҬ��*���:�7�ѣu���,��`� ��[��ƾ�@��8�u{��vK[[yd~Q�z(�����N�VX9�q���G�yC�<�9���Ou�@�����z*y)cJ�z�?����&��(���t�K�4�coڜ�Cw��/0�ÆM�/�t�~��Dq��.+�X��d�	���~3<�53HB,�L_&S[����,ә���+O��J�1���[�W
�.�[d1̐���Tў��m?�	uA�y�K��"&RBF�Z�rA�e��s��(/M�$�MPD� �'!U��惏��8�=�=���M<�I��S���<�J�������!����ۮ���<�n,u~;n5SM�>��O�B��0�S�؍.&�m���-�^����ԍ8i�>ǋL���u�6q�#���_�	����M��ؐZ`a&�"�/���\}��Ƃ�c�TfA���Yڻt�
Oe�%�M��Fv�k���s���_�]��:�/=�:}�L�z�\0S�ɯk�,���=F� ��b�ZW���$ހ �m����M,�������YfR<�F"SH�3Z�Y�b7:;'V���U�o2}�k���hp�"���X�j�t)׿�����m�W��m�q�oJ%��OqVzA�Ah������S��x
�c�4��x6��\�%����'��|I���m݄?�A_;dX�F�:�ŌA4� @�ue� ���Jg��m<��Ϳ{3~	�X��sH�(��A&����D�C�x����!4! �Be9
���s��M���q�sŅ���~��匋\dȬT�v��3�@�ߏ�,����7Ч�zp� ������뀲t�P����H��D֊,���o�G<�"�I�&�j�W����n?Z!9PnAq�8�*�兀t6w����U_SC���D��p�ܔ�aȎ���H�|�B%�9��r!���3`V_tJ�����5A�#�P��j}���֧�O1E�p::�FkK~ut`G�>�"��B.��G�f�	T�����4A6�j�����.Ns	0ʎ}�e�����Y��a�5ȇK���v@^g��޼���hh�TS=+
;:3Jg��Qs@�U	n2$-���"�d%�"��N�b|�s��t�l�͑�T!RVrm��3:��_�^o� +����vx�r���}�R��0�@�L3�oA`�}.�*��تz�Kd.�q����C�:;�l��gFR����B���Jl`�p�?;��9�� �`�������R����s9I�5������5�T���'vI��M8�;����ɞ���D�q<��4�	N��Yt�k�1�b�Q��2����z�tĞCh~#���
]ɞ5���Y���$�S��α��n,bR-��h����M1���=[ߚ�����~��v�$����wtu"�To���z6���>�3��5lB�Ԉ*!nC;>�V(Vv����eQf_c�h/Ǡ�!����vBV\A~5#�zΑ�_J޸q���խΞN�\���h����a:g4S�֘	
Ee�W�ᾥ�%�F�[d����Y[�G���	3��7��C'[YX��{L��
͊|�Dzu����J>��c�;�M��E����]w.#ɘ�b�����(��v��]�d]�>T��:��)"�+�b��U��-�pǨ�:����p�#�{�)A�ms���>q�ڃ���Qv�����NÔ,K