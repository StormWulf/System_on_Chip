XlxV64EB    3b0f     f00��n�`IJ����\��i�%y�/9��В�G)��T�6Y��@䘈��;_�\��g*���O��]������u�sG��ϳ{"��\u`wۨB������4��>;s�G� �aӶbvu��|$*7�?WjA�R�Ʒi�Y_�WD���o��,�aZG�և�P�݀�z@���E�����3`:����t��Ke�Y�d�����|8�Ac��3|i�_q#'����i���o���ߜL���?����� ��>9KЅ<cw�|��;�kb�UA@}�N�'K0CcB���I��	��N��%���?dB�o���ê8cdۍwB��t��5dY�}d�P��۲*�����:d��,W:m��ڵ7�d��1��6�Rp�|����6�����e�rK�鮎�����	�1ծ��f^HJu�gD�<��M�Y�c�΁]��*9�_��}D�H�f̽�5������.�wiΒ3�ؕJ靝�u�օ�����.�� ���t?�lH"�ĸ<�;�/oRQ�S�z��1���'7u�4�r��fC�� G��XncEKǔ�Y쑯�鮴�@vVُ��<���d�Χt��jI���g�����0�c��pQ��������$��6/�/7��kS/nK�u��5���܃P
)ts�%��gS�i&e|�w�O|������1��kQ+��HA����Rt T%��.ƥ��F�A�?E���B�a
�<�+���
x�SA�ŗ�L��|��u�0?kj�ߥg�!Pg��"d���}�B{H�\1�H$��zᡬt���ڕ˛��z�V���lϾ?*��}��ť�ٮ
�n6���Yғi��|��~k���H���g���.%J����n<q �j6\��P5��'�a����[-���ʐ�{g�8����\�N�����0N�H���"�s��@1a~�?�N�Oe_[P���r�W
�_�;y�7��o�WH��� �.�6e�݇������]e�T��C�v(\��;"�+)��׼�P��`m�R)B�4ȁ������� �Z;ڻ�U��>74�}N�7�S���t/뗲�	�M�"/���$vC*� ��u1�rx�Ʋ����5ɑ��44�����},N4��QN?k�g�>鎖Ul�k���:���pnU{����|$��7|��"N�]:���t��@r�5�ԲmԢ
�Ĥ�$CV�(��w��y I�~ >k���o%��^���b��Ի�.� R�)�6�tu�0`�{+Bڟ>��'�xx����D�J0�e��y����-;.M��ќop���_&���"�l* �$���8��A3|f`r�`'3�փ��Ѻ���Ŭb����Cv��'�K�OP��q�2bq@����?�3��u������w���a�Ҕbq�]x0�ѕ�1d�ؒ���`�������YnuH!$�0}���I�#G�.̅|o�~_��~\֍f�OR�)���zŚ�4y��V8qol�B�ρ��R���&�_F�<�]�T>9��Z�N���{�����:�p:c`(0��~ۥ���A�g`Ԏ5���w��>ZzJ�H"*�L�@=�)�C�z2 ����N���Z`�n?��#���H�)k|���*���]Ѥ�R;�M>��2~��B��Z�)�ѐ�Q�֍���O�Zc��r"Ei^��q&)��jލ`����N����(!T=�g�45�P��62��Qg�ɱ6sl���6n����~bϫ�	�N�r��8�E��F�=��]��0��!�IaY�!}s��Z\d�w��~��W�F~�6w�c��w���إ,�hA�E{;��l/H���?�b|��٣2_�r�3��!��
e��b
�}��y.n`]�#�� �O�|�	%�nj��q��ԫ"������2ՠ�p��¾�O�ν�]����*f�	�4x�?�e�ͫ�}�4t�QN�	������^���Ct�J-�?�!�L�a.��Y�W���f��#�H�ϯpedp�\0z�-7tV��xH��;�sj���d����_���nঠ��RH=��]0mw9`}o�P�T����A3�F
��m P�်\���Z���� cJ��?��;��M�6��s�v��[3ȿ	Sq)��'
����IS��O�D���y�t�:lJK^y�~�X��x�_:?�v*�(��Yj�>�UX�h=�m=]�iЈ.�0��g�MQ#n�`S��� ^�2a��Ôi����o��*���g`��U�f�J�H�!�m�Qz)��di/{}WʅE?Dc�ӿ�c�$�Y�1	��!9��5�c��J����\��:��+g�¾a�$���|��	�S�-Pt2��EN�Oo�Z�(�,��1�����kH�'&���j%�{�k1�Q4��g��]����<����w&�P�5�
e�4��3��T�HI&L¹��b�=��asǖ���=��X��!^�'2�ʃCS	����C�D���/RQu�}?�$�D�Zb��_8�c�*�� ������i��6�����P�3���e���#��Ji�yyb��0��_N�G�l�Au �O���z4<�᧍�a� ������o���c*!��x�,�1�w�s-`��X}5l����� ��IRXGI�N��|�Mln2�������7f$�- �9���j|�|������B����� ܆�%����O0M�lX�#0?ؽ�Ł>N�����Me�Zў{o4<�O��}ceYF�p{����q$5=�eUz�Ɛ���Y�پn�J�����t/4��T��<sn��|^�n�����W|�vjq>FC�2�"ҥ�`-����3�l���ZT("�pB�f�.��ކ�����hbmv�RJ��'(��0M��<����Y���nťc`�m�\�b����:�";s΢-��R�XcG���:��g�S
W�5X���8o '�=��O�"�y�m�z�:*����xF9!6�.aͣB`�ې�2Őm�4U���{��!�P+��ٰq��<!~1��g���8,j
@�H�;ѐz��� ��"Q
�����H��r�
����?K�ɝ�$c�M]�����Gt���_,Q�>������P�7��� ����	t��V��렭W�#*��qߏ�'T���o����]~+餳�62����h���)5l�<g�W��F�g���~\�oCP�EN2?H����*�+A!t���7�6gn�Rty����KJ[Z��]�g��65^Ԫgk��;�W���7���?��{G��� q��dҩ$����J���ɣd��h(?Nu��/�GAr�@V�b��?�s����Ry0��hm��V�D�6��B���㦌�f�mƳ�4͡?�v��&"<�T�u���/�Q5`{��j�T.C��^����y�<�h�7��G]�~Z��Q��u�=�G���q��>��Q���zp ݐr�IR>ϧ�Te���-�YW؝Kw�����Tף\vJ�@��' b�R=~�~�K�THF]yR�:�����A"��Y�|zÔ?];"%%�+D0zej]D�C!��xG�%��w��Z�<�px�B9�[��;ymt�X�J�Eɞ�kĀhd��:�rAa1,�R�.G-���C6���B���W�2~�y�j��@��jS�M�d����<gCd6��(^��5�$�,=�)����N�p`�)�5����q¼k����Z�z��Į���Ζ�z�.���XR: )[��+��(1�rsY5a$��D�ּ�k�j$^����^��