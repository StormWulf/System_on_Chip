XlxV64EB    53dd    1130<l��6�w��e^�EX�����w��|�4�O1�h��2�W	����tUg<�ٲa7��Rm1�M�6�楆��q���,cم #!KW�x`4V��w����Z,*7�i�\$�����gŬbW�B2>/���+���}RBќ[��?�J�����c�@8��tOϩ�6��҈�ϻĀ�MN�3T��,z�t����|+�`o?�MW�?<o)�0IW���z������i"���=���;*�y��ֲ��Ͼ\'�d�J:�X�&y�ѥ�))�����d���&�����4�%�m�ި�	N�q-�)��1^_��)oroŮo1�NW��؝�ݪ_�����>�����ʽ��V�9�~�>ҡ�5V$��s�t�M�d!�-�C�����%\#R2�B�2�gMfP*����^t������u�cj%q� �|&{���	^`!#6��Z!��ސ������+*S����f9ϗ]��y�-+/�J���e�E�w]������ۉ��mnk���XDc�))Ȑ^D�O}3��)������0��E�6��<p�]���F�6�Jً�,�ᮝȱXIˇ�8"��j�1<�[n�	���3�_n��|�E��a���`��_&:�')�nh��ևk�[r��K���˔�x�ڬ
s��8Z���5�@W��⼸�j��w[��22�J���'�=D�+6<}�J@��6� �.���*4�@��k�����I}
�e0�ߵ�õ=]<\��Lh;����F)����Fg�;��;_�O}�]�6:t��\�V݉�X��f��]������Q-� ��/_<l,`D!�����aʈ������E^�@�ɉPt��Dtg�e �����.�QIلnfQ�گ$lOc�c#a�y�k�r>�	�b�ؒ F�
������8'j���r<BTec�'^��i'�l�]�^W�;�5~��"�?�S�l��|ﳇ��-I2�
n��3�1�Wc^O���m�W�S	��,��=~Z��D�l�8��X)d&�G��>�qof��1����?ӬZ�fզoǕ�$~�-KC&S��:f�vȬ�\�6�èdo.A�`�1C����p��2���k�Z�-!���Y�W�U�8bطi�&`Q��� �^���!Z���mN���
�?2ϙ�7O���� �,Hkr�ҹӻ$��m~sV�q�2�C5��oL���D�~\�dHӫZ�,ҡv���""��CϬ�u�Ŏ-Uj�
/O|��=s8�j�����Й���*� </&��g�9�T����s�$Ǆ�M`�Ӱ3��n��)�����_�Z�+v�㤱!a?Y�n�}��C�Oaa�4��?C���~��6��c@���R�aAS���I���q��:(���)�����Z:B�2>d7>\J\�Xq��y8�o�s��dD��'PB�jd1e��_�A�}Јd�A�KXu2����%�aYB>��t��e�?��rA�����Lsևf�x�����X 0�Y/EZƄ$�����w=vMz!P��Q7'18)o���t��1�J����]�I�?����L���{O5�����^�]�ނ�_s�A�0�eNP�Tʡfš�=�9�eD˺���rl;��%jTN�.��Q���X��ξG���iϳ�ϵ�Ҝ��sGW����E��*�{����h�U�,�1�C<���6g�eE[���_�p���
�>l��ෝhH$�T@�Q+���qAa/��/�h7����7��)�C�s��Ew �Z\,�F�S Sa��v艧*���֨���uA
i=|����F<��m.����5+_�Tk���8�Ί�m(� R�v���bę-n����m���Yo�LWV��M�M�qH1�-qۄ����z����g����:R��&�x쩰��O�-��٘���˟�BlX�?`
$�l�sڢ�U�fg��-�d��8��s�R�k�n� l��I�y[�u�Lg�hX��y]��x��9�j x0�3���6�W�~��@��p���s��`����E��i	��c��~{�עXu��nKi�8��?��~e�2t��Jm!>��K[��7Ԁ�&�*5	�A6]�}q;x�)v�
L%��h3y�D;�}���zc�rdZ����vR�vĤ|�ml���9f���� b�������3x�6�4���g͝����- ����V���ZĎ�ߪ.���1��wA_RhOB#��Q��N�_������~'n��m�V�>62�F}��y�򟫑v��Ck����T*��H��D9-šu#+�iq. V�E������rI����a�%��+*(Q��V���ZU��.0��6u��S��Q�^)߻���"!DE��+�85�\�*�8�Al#Z�(����N
�����5��"�3v�C0�~����#k��[��L�Q^��I��¡����閭FލW�",U�����n%�O���0��S-�~�m�Kv��g$�/.|t�f�0N�V)��
�$�|��b))SU����6�j�"�^Ӡ�hW���~�Cs�o:�3�A�7[�e���Ú�J{-�s[a��e7t'�b���Kc��ERc� �i��=;;�|��9�5�v���#��5���F��ӱ��;P�5��\D+��=���£�[ag�ؠB�w˪�zf�'�_
�ށhF l�4u��#���XՅ����7����b2Ƒ2�K��[B8Ys���1�I���2��¹�qrYn޵q~kY���@��U�mW���ꎥ�(��h�=��aJ6�v���� I�}aLp�kCE~>����f��RԖ?K�_��#��xd%�06�$���[$��SCf���PR-t��{�+wˈ��A���b�Ǡ��H�T��.i�6i�o��b��/J!��sFGݎ��U@Z�H%H 6:T0Φ�Nt6}mІLF�1�W����opq��h��4w�'�Q6T��	�z���/"E��:�Ncg���ɬ�	�����OxO�x����ϛ�Jfjч�D���ī�6�l��@ ��Ġb��bv"��F����sዀ���jw�3*.���*Ӭ-����by�ƪ��Aۢ*���fG}����\������|�K��,�*�ۑ�w��\�q�GV�B������a�)(t����g|"�u`�<!͉�^����	�#���W�d����d�D�;�d+�Mo��WE%. ��v�k�&�wC�u�4p��r�<C�i����6_�r� B���@p�Y2e�	�q��ħ��������*:4	Q{���(?�Pbl����lwp�'0��5��C��i�f=sG�JK�C�l�g���~���p�䘳���G�? =׍�?��L��k;�h��'a��'�s����`��>~�J��[�4c�2�ڣ�ɣ��g����."�"���@õV���#,�yl��@�ǀ( 𗜉�X<���O�#��'����:�Σ�=缱_S���yy%���.�&�/w4��������K�ɀ���E�u�V�FF�o�d�ܯ����&�{�H	�!Q�����ӛ�&��f[u&�f��4U� ���>]�@��GZ��(V=�#�H�]���R���%#v�5�n��8_	$��WF��q�}�Qu��Ȝ�P���v��ax4j?|��s4��;�R�8���7�T4UG�wx&Z( wl��t[���H��x��4��p�E�8�uL�3�A��=����l�A��.��韋а�����j�Sy�la�c�n���2r�y����{cD���
���<��Tp}a�	KT������fo��]J ֵ>�+�\S~�k��[xM_��ׅ05.�O�ʮ�tx1��i����m�Ȯ�f<2�'��I�5Nޖ�)��hz�8g�)���j�nW��[���k$�(��	e�� ����+I�CZ�;��-����?�=bR|S���gkݪF��=)t�࢞��	���x8��Lp�) 0�v��ޡ���^����_!��/��p�A�wP�Pҡ��CZg��qr�i�����2����}[�˱����!`/��udԖK�\q�{�H_�^��h�6e)�/x��\b�>a���F�{W�>דD��%c�G����L��a%����H�C%f��f���!��1�D��Ά�)a�@�Jo%��QIM��|��^��!b���H��g�~��-�L���ަ�lyة��Q��ώ��f\� �P?�ȉD�銮t��2��G�4�����V�!R-�}|�z;G��=�ht]����ZQR���������ڥ���;	n�ӗ��yܿË#0*�?�xRb���f	��]