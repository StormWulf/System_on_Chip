XlxV64EB    fa00    2ea0Z����y���b��K��i��#N��R�q�["`VV���=`@�b��#I.!�
N��Z&T�'$���5����"����@���aԩ�LF߳1w�P�F�m�n���j|�-ߗ3P��]<�w���������V���48�@�JBؽ�v�R�ƹ�Ύb�C�5� t�=�x��^��Ub�r���ݒ{�}��b9�}Q�Zc�������1� �L��T����b޷���mk#T�\��Y�>�����.]�D@?�����������O�_��z��{\ꀐܛM�X,����8:} ��<�4��Kd�M���z_�`������Wޞ�׭���H�k"������3�/���M��+��"�·�p�ȸ������m�!�l����8>��[c����ɛFrB����uy#'��!�����v%t�G�
Uu����*�v��Ě(�u@��\o���o����v�@G����ld&�����[�8OnLQ����lw�O��0d��O��(���Ye��y�\����h��
3�?bJ�OM%:(�$�{��/�C�1f\�&(8���b�n�	��ch.�$nUv)�`��`M��6B�A	����UZ�<��|Z�-��W���ҫ�tq�n"+�%"���&���ٗ�Z	�w��n��@�Vr��Ѯ�#o��j��"��gK���Ht�Wn��ݙeB���Ǉ�:4�#�%��vҟqWL:`c�x�RݟYƛ��E�>�����Iwjk�J�B���ά;K�gv�"9*4�k��=��҇�nB�g֠d߅
�e�-�59]�y%���`�u�PYnl��̣ ��e�3P�����?ɸ�	��i���}p�|� O~���~vyVA|��v�RZ�	İ	��.��e�2�Q�@�~Z}�\wvS^S�p~ˡv�З�Q�ecS�pԦ �q&�'�=��2w+��f��͙�c�������.
%�N>M��B�K�JXqxv��EL4Z�gOyMb`Еِ�/ȫX��:֡d[(�[��f����拡�Ubi��"d�C���"ןNB��7�.{f��̊U�'V8n��~U��4�~ӆ��N �����tP�Igci�T�U+*G�*-���{ ^���!ִ5��x$e����J�4-#����i��-���~��UP�"�P�~�i�v�]���f��K�o���,��!B����L7v����k��O��I%��s)���1D'�h��5Uin����ydd4�е�-���&�gR�����������-�ڋ���: �r���̤�V�
#�j��ƃKh�t�ב?�����ό{�s�Ѝ� :�9��/��K��b����Zib�nZ���;��%4RC)�[h�w>����O�l_4 ��!�pW�2�ʌ��Ld��T��f����6r��,t��X\D�h_�j���_���=��3��!/pt�#��rx�B/��*� JȰ�
���<���q��m뚶Q��g���m-�ڣ��̖[�]h�-���D�2Y�k[=��i���/1(@R����#J/��c�\�A�K�q%��	�ɥ4�U�6��AEY���\TQ �h�Dyf=�Q5p���Z�>4t��(�3pֻ��Ɩ�}��02o6
�I�~�C�&�T�N�J����ۋ&�~	�4�<^l��d�����}D/+ioZg";�]	�0���	.�`%���e"�]��[+^��a�/��{E�\�+�e)�*��os�� 0l�
�����v�P$���tT�����O
<�G�Fi�|�hWo��pB���/*ʛ(b-x�໿�ʃ$����E���K	ۭy\����	�b�dp`��Z���Q{3#��x��Z����t��'J���C����c�/pls��lL��H�k{�Kg���Lb��C>Ƣ����瞲��(��
��֏4�\�$�n�!����gث�mT*�Y7�U��v-��:�v�0�K��c;��B�.�)b�%Lט���R���L��N՘�Y���WV��7�DAn�$��]<����B���z< �� L�т����R>%w��:��#P�,5s��1�3z� 𵸗*;7Զ���|g�N\~����s++�c����mG]���ԏ4k^�+��y-l���>D�s�0t#���c�������6�O>	�P���,��l���l��Ej+�Bg�K ;KM�`��H�,:-�Q0hUc���qv�CXW��ز�T�nM	v���;N����Yy�a���H�V}׮����l�j�Q=�p)d��:b#�l0P δ_U��X$Q��R�A��4�{������ w�#cwԝ�~�Y�,��o��I�'g8߉��jps�)�ğ2SmO�383V�vV��L�<W�,(m�VD����33P�K�AP�DEl��+�_����q�����W��J2ĸ��A�_Ģ,Y�XV�9���L5f��<'�K��~������SS$\j�bwG����U�r�mb�5�T�O&0��u�-"�^~r��2�B@a��r��بq%�|�CFu���B�w�5��4���>���*�^����HI���D��C�pʚ?�8h���#l��Hb�C�X��5x����
x6Ii5�6���_�d����,y]�� Uq�H����߽ː����RF>�Ak�ۏ��@a����d-
��A,����>�I�����@Qv����g���J�: �דᤢ����q����f_��ʿ���Z�*�yY��~�9r����n����Lx�S1��Rv�5�c�S+�3��]U4>�����4���h�ƕ��g�T&�D�-��Iw����a���:gq{p7j r[��.��GЦHX94����󵰞a9�C�\;��bwq?BS;qp��;�TR��ۥ�*`�
�i:찈���=5t��6D����>�%��h;T"q-��&\:��f vy��ʆ�f�9p�y\<�^s�Z>C��E�5Z'��sIi��}���Ű���T��0�#<�|������j"Ѫ�����:@O��S�I�[�'Qa�VƖ��dbaf��mٟ���9-]�_3y��,%�n��,�qg��⑞{�ޟ�D�4۾_U�]{��E� 3	�@m0܂�F
r�jtѡ*M��Cx���.AG	B7��7�/S��\,EE�	��bn�}�`���������ȮM�j3/Й�S��dd�
*���q�+�<��h�+�1kޕ�|{�V�J��Bv�;�w.� ��	LrK���8�X_��Y9孧��[+�jd�4Kknz"�IS�LGAŤ���xrNy=�]k�T�q%h�sw��{�Y~>m����pI�O�8��r')�;�8�N9kF_�jE�,�:O��S�]�iC)�?��4�*�s�f3}���'.���mEZTڳoƶހ7��67�����xȗ��q���ʐ�F���m�1FQS�x�	 i����ҝ��ih�+'�Xb�X�Xn~:肯�Tm���Me�:�Z�u0>�� |�0�"S�*��|�\-�Nh��v�p���34�W��I������8%�z�z, ���6��<��R@�
i��D6=vv�+����s*Xa^}^N^�EL�4ь:h�I����AϘ�M���n"�`#��݆�_΢�;�Z�B�ȏ>}Qqf�ȗP�	Ptn8�}�H>aP;��1o��l�R�=-HF#�*��
[_ז�ӂ=AFt�N�Y>n����aE�������8��C7��{='�Zu6�U?�h���e��4�t̜��0W3ۈ�'$@�J<�*�K��:*�8��rU��{�yۻ�WR*�r�
���7Ok�1/yL�#7��u'����eJ���c������O�����00�x��ڄ��-��>�����ø�����|���'*Z&��WR��rc-�j�L׏�'\���h�C�_���8��ポc�<�1u_�V�/�@qp���)�W��`(
���=j_�/��@a�%�R��kH��7��pHP��JMy�|���H0���؏�t�!* bMm _�����sW�.ϼ���!<�_=�b�MNVf�=���Lݭ�9y���`��?�Ca�J��q����9�q�WO� sM��ԑ�28���l��Q�H[�t�1LS�
����n�u��h")Պ8+�&A��	䖮�_�\��������]�e�h/��/v�>iC�N��X���;-����F?B�����P�T�h��J5�Jc� Ax�'�	JV�_�L����́�ȫ$�d�yў�C�.4�A����g>����3I��3�U������y��G�� F�����U����/!!k?M޴�9�>a�-<�Q4T����e���o���%�h�$���+5����R�񆇼F��
zQ�]9�?������I\�SG	7Is\� W����C��!�Q�0��]�c�I�g�E�c�J�X�uZ���eQ ��g&b�*k�7N%�s����R��U�a���]V��_�N.;���nZ��D��x���M���dJ�b���������G����>T5mW��g)knשu�U^�������o��r�+P��<���[���H!`,� ��g������1�Ѻ���= mZ.�=P�q$&K�u�|����+E8N�ٓj���QzM��F�t1�T]U��&"j����f�C�!n��eq�K>QL�#�_�V@Ze ��]')���y�Noؗ�T�zv]�U��-�Yg9�_Oω ���%N8vp����hl+glAwr��m�n�_�d�E�1�q�KG��U����ԁ4ܮ��G��tS!s�G���k��;z��S� r���{t�{0gw�Ϥt{ҧP�3���_7�mD<�=��|�0��Hتc�!7l�R�ŭn�b{(�c@�6D�M�)�I^�c��Տ������z��7t(���o���	EG��|�����~Ĵ=�R��S]+3;4�dm3݌�⑁�B]�s%�0tm��`���Rj���D�s���X�b��V��5�W��M��5�N�q�,�C�
���qKu�/s:���|�k��0d�vZ7�9��x��E�SL+����$7��V謁��P�5vΟ
f��v�Μ�GP����/���7^�V�����������A���w��GP�� ����W��%޾�P���d����'߽{i��rQ�P�󄕨l	�}sO�.��{]�M�͔�&'�]ZY$#�����=�%v�n�ኮ//2��ix%����5㐧p�J�s�T�#i�h�Eݰ�l�Z<$�ӢO�����H4	c9�}�`��ݍg�W�@����L�<���h���"E��$O��:z��d��naa�����SXG����~���C'�Ea�$z�d�'�E������{ޙ��uz��R�F������D5���P�] �	�y��ÿ�9:��~�H�]i\C6���46�,r���I6��C�x _��W}K��w�)��������zE+a�բ��	d������e��yUV�M�m�UV��g��C%�蹾,�:|\��#��-3���?�2����yv������ΐ����{��K�+�j�@����3e8~e���c����QRIֈ�!�.W��D�6�r�sj�,��<�4�9��e��5<��Q���\�����ӌ�Ԋz�����y[��0�P�w�aF�pELoW좖$�V�S���� b�Y/��SYkPr�����-*?|C_����]9�2ե䳪�g����2��> K�4P�;Z�@�Qڙ<�@�K�����MH�*�0��-�����7��L�^����&���vE��?�~���gs����/�a8�����F^������+���$�R���'x��d���%$�	ƾ�����2����/�v��#�Ԣ�dya��^��Y-�{�w?Q��<�v嗾,����(��0�|�i�;Ci��c��9�#��r �8�)��+�T���c��=2��s���yj�� ���Σ>^f���}DS��h�9Fve���*bȀo����2|���VyG!42�lWA�L�i�SȰ8O������C%���z>
�ڤ��:����wvN���.��i��Eq��<UԚ��3Lu�V�������w%KEMȎ z^���e��9K�D���*_WwĶ
�sn>�!��"�]W�&J`��8�*e��c ��~���LC����!{��@|J�,Hd�ӊ�+Z�z��r��a{b4�6�8u�0���'�"yn4ڔg=���m�#�}$�����ꔿ�Z�];w��eM��S^���xgT�/�����<�<{�m��^]״������<�D���G�&�6�y���s��Ԥ��9)en9Ѡ�Z�>@��Y�:�
����CE
����K�6���� �.7nW�w�͈
r�}�ɒ�.�h r�R�Md�Wvu��v����u#�2���U�9�65}�K U0��~õ���
�OF�������0
�J�*��O��7�����,ϔ��Mҙ���.RO���rO�lR
{��α������� �#�w22��u��3Z�qXͨ�1�t�.zHS��{� �)�J���:]�``9��w�%�&�ѷDm���L{"&��͛|:���Js�Nm�K�3FP�hk�f�5A�B;:��T� ����:�hn�G0�R�@��'O���|���*����S�e wy��������i�z�p�n̸�ej�e�Ԏ�_nzs;��}J�"�$�%�~\���'�J�$t�m�d"=� 9�Oujk1�D3y��m�/����?6��6�\��)2Jv����>�~�f�x�{M��ߧ��pi�3�� ^~X���Ȼ�����l�����I��B3��m/���Mr�R��z�4f��pb^���{X>TB�P�^�D����4��A�B��Y�k�jJ�-h��zh�C"c�u�"��
���K���AA/��NSV�+��@צ���ё���:�|@�g�[��Cl�?��\��G2�į�5Ȝz#՚��0'�ׇwq��!&�/s����Kq��->l��J���&��R��9S�\��C�/mu4P�����vB�r��D1���9j��G��,cӇ*�i��~O,7q�����	2��lčP�3��3�O��;Λ�k�P+E#�n_��(P�4|���^�**0g����,�}�ԙ| ���/���N-���K"q�����`c���@@#��r:�+��%U��	����'�'�ġ��
H�� �h~g�=y�=��s�N(���Z�yP�[�v����
췪��.i�1���'�3%�	���`s=:va\��o����Տ�j0�j�,�8�p�����+�&�^��t��F�����~v��ײl��:x6�� ?�*nJa�&��bGS�(��Y�h�!` �+���o�����%�~�F��iq񡶬�S�Z4��U@,�w�X��?�R	@�
5��8-���u	��a���`R�e���[�1<�:�?T�J$��il=m�5r��L����u?e�PM�
����.�=��R��ga�f3^��=�4�l���~2�>z��"ŧ��i4
�]�7��%q���K���1]��5��p�oU+3�� �Y��й#��9��5Xn���F�萡6@�3���YƊ��1�5��
�(� �¼{����A��Y��1+Uۓ~:�nE�f��{���1�,�����M�h���@��Y�:n�DM#��\쉉]߃'� �j�v'p�xm:#���w��ȡT@׋STe�����mP���x�G��t��_Z��] ��G,�4ID���S+�e
��h������L<9f;\����jm2xf����;*=Է�p�r#0��kR`o�2�o4fǀ��,�DM�6}_���թ3�o�mjT,H��h��
���5�>�y}t�
��.=E@I�ö��9���������>�R��c�)*r�jŮ���o�a-$ߡ.%Ez^����Yk��!�H����D7=;�q�^>��@�}� �x��Jx��qȨ�_���j4�>\:+r�Գ8aM�eb��(J�)��2>��J�P+z1����+^�S����՛�l�ٛ������7�C^EOZ��'��N⟜7�!b��N�Ã`<Z �l�ɐM��v+=���˦�ʏ~�����wZ�X���5��|��`�<��)�[Y 3G���-Z(uyX���5݇n©�@�An�M�����*Jr�1<�Y�z������J����� ��}�!�FMɋ��7	-M�A�"�5e��Z���\M���s�WA�#��v��F����T�AG5;Sv&��E�[��b�g4/�V�t�v�>��QK�^����Y��O�򰆴���~m�O7��;i�'�!��;��O6�?��^�b�5��_���Ŷ�ˣ��w�0X�S��2�"���P�gU�Y�4:�C���/�L$,�^��&\8��h�I�oo.�^y ��Zg�cW�uF�o���|-��]8��&�i@g],�.���o�$L{w���z�-�����-�� %���Z�`��;$��5�]��5w�.R,�C���QJ��BM����\�V������sL�ΐȺ<}[������̆n/��憿'U~7H|��D�kr��;�h�-�7�鱾mX/�=��I$�d�π��R`6�O��r󫾇�>���\%�2 ��$�J#��T���9ud��Ka��+3�j��WuF86:9vv �:��Iu�� ��]����r�{cY�A�Uh����8�NZ�y�+b=�%k�윇������H��z�w�j|���%).�����l���\�v��~��%���=] Zr�[xv�W�ׄU�A��=jLSw��рt<�gK�x!��T��%6f�I��c����$�p�pE�D��R������n�$�䬷?D�-R�t��ֻՠa������N�Wh�8g����m,�N�ʼ��TU��J���hF]3��L��G�4�i�0���L��-�Ib����]M��ħ,I�[�j��K��|R>��񒞉钅s�M `��I�9��N�l���Z;q@�SC\���d�f\ɦ/Uam����eohA�ʫ�e�流�ZIZ���^P0<#GB ���I��$����ӻt}� �U<�*�F�a0S����Q��?7��/}����HJR�l5���<.��Hl��d":�m����2>�2�@�*uy�9�3�^��Wّ��'����A��
D�[t��V{�]#�L�(p1�(���Y\�ۤ	�V֎� ����,~���
�J����GN���Y�D����*^p�ͨ��x�c���Y��Ce<���H��jX~?�V^7�	Q^��[n�q�Tuu]�Ϙf�"�oq��@�G�F�H��KsUٝD�?�z��J�RFk3������|C����	�d�M��-�W����<p����5nQ5=w��?\�W�V��{��0E�5�a��m�?�m�*[Ǉ\Q�9���'�z
�p��DF��&Z�D̓��)��|��*H؃��H�Aq��+<����#J~���{
��ߚ��W����V�d����f���;l;�t>1�����f��|E��Q]X��]���p��wz�}���^ĸî�ؘ*+���Q@w��N�l�p��0��2\��X�A�1nA�B���q]�:�IT��&� �J
����ᏲHb$���u�U-2�H��0n&|K��dgw��#��sD��`:����n򐊾��U�*�։�Zv�	I�_��W>�f@�E��䩡6_)p�	B�n͟��fe5Z�r�^m���Y�l�!̨L��2hD��lI����H&-��b/��4>r^o�!�OӬ�4�L�X�GڝF��ÜPb:/vV������J��D,p��PB���<�e�yf�J
������=�C`͈b�����H���˂�>nUꞤ�Ӎ�$��j��cȻs\:�IC�|�O��	Gz���P�YmѨކ�`6�<
u���3�����
ځ	�-
e����}��)�кL+Qժ9�u>k��~��^E��&� �|�6����NT�6���ңv�[��擇%ޖ1L[$��Y<]�hȏzi�eq2:��](��B��>:U�:�~�8�9Y}�@TmR[ǜ�`w8�4��[7�Y��^�%� �f�G)7֫�%���$!(�rE����!�ƻ�)jN�U\*	D�I�3��.j�̈p벉 �F�a?���B͐�0�I Nyxu�0������(���ĚYH�"����4��B�˅�l��e��`��^lP0,�{��?umc5�`hu���"4������ٽ6��[{��O9QUG���{���]�n-Ns�\) ��CW�<���54�o'"N������7*FByJL��r�/Ԃ��(rrPW��{��u�5����w68/�lJ~n�텍g+ ��2Ւ�rcħ�Xzf ��K[�E����;�c������i�N�z=�zI^"v W�>K���Az�'
�=?��<��=��-i)��{�d�.�7_
ҕ�Fman�o�C�_pQ1h��L
lliub�X�~2��u���L��3��	�!"ᝉKZo\����C�z�7�A�U��63�g����sVw-Q%��k>�ϓ����4�?��(�U�=QԼ/�1��
�"���ܖHj���"2<e[̜*@��{Φ�v�]�ю���]C�QI��i>r[��c���@6��8��C�:lC1�(u85Dc����k�vmQLI�Ϝ��N9�e50���G฼AmO2Ų��9$�a�z)�-��Ry�"�D��
���J���T�VQ�8?�
��~0��4H#fd��S ��l_t�׳���^s�JJ�v������v'Χȳ�oJBAi&��p�-$pr*@D�Y�o�=�����a��ע��nX_}y�@͟���Y��أ�!���*m�Z��b�w0/,����`��d���D�����|R�x��/Y��a<��7�k�X��������2�خJKk½⌰�<��
0����BK���d��3�v�zyK/y���7:&(��+o�x��<�\q��Ô媾�B۰Dm6�S�yvOIW'U)^#�T5�2/���`t��k�V�x�ى��������*:P����Ȩ�NV�.;a!�����p��e�x���y��_U�v�S7�F!R.�m��Hb���Q���D?ܱ�+�v�ƶ(� n?��"�l1�#��� �V�D��l��/Pd�5�n� ۆۤפ�f �l��y|��Fc��^�әa�!����@���A3~���N8�����n&6����B�;��EA"�Y����D���pS�o����&�T�z�D:����ć�����ILy|��g�L8����d��q����ky��,��ӷ�lB)b�䥹+�U,¯6j�^D��Y�.S#��H��_�5�^D�#Q��Ɓ#s�=�C@�	�N"��x6�+q.�G�(.颇0��)����R�K�%��m<QF����q�K��-�����3�`Scj/�F�l>�<�g3�~j��8�|.��{�s���I!S�oT�f��l�RXqi����#KH��~dW�f`O�*9w'��"�q��� �ItRTGm�Շ���rc�F��lX�)����ncr�M��|�	4r�TTj<|�Z���0bcXlxV64EB    fa00    2bd0W��Z:���{Tרȳ�s��u�p��G��u�]��}F�f`��F*�
{����@8`保���!���r�6��'��������:��T��*m�TtO��`�>,L����PP��6�*�,������FPD�q�-_९o�~#嬓�ksA�zm��P����u4cKa-�*�Ӯ{��$��ٷ�3�T�r��uŮ�ۦ�K�w 埁stC�r]���9�ޙ�Y�1H����K�?�,l�[�;�ܥ�6{U�B׮3g�%d��uWwJ�L�Y������-C���+��0��x`�R3�|���P��������H�g�s�scڹ|��(���$����v&���]�ڥ<|��!����I���b)�=h�g�a���騿�A�t�M(L4b�� ĩ��睫'�h��ߐ��H&>ڻ'��s�U���]c����"�7���~�����I<L;���w��ڰ�H�\��z��VA~�z7��
���o�N&�S���<���D�0�s���B�̓�&UzBzUNP+)�	=�μ�0¾�`�j���)@ 5�Jx���aeCԦ�
J7��4��F%�-l_I���<��aL�Z[���{��`�C�j���
6�}YV��@q���qk���B�n�yi���b���M��>��n���tW@���ݮ"�hPG-�\�\��2Q��^�~�Oл��_�\6��)���=;�Ԩ��3�Q�
��OQ��4(�4u�B�V�V�Q1n���\�h����]h�>�G�����;�x�f��~�F��},�U�&�T
��Xhڏ�O���W��|�\͛�7��� $����7|��y]"��l�ʱZ�c��G���	�$#��V�2�8�Us���r9��\�a�TU��'�y���Ө>���Õ���ܾrU��G�7���f/$�\�E��h��X ��b.Z��MP���D,��Jyx�?��Z�	��k<a9k�庌Ѹ�r���)�?��*%#T����w����K�]t����� $�Kʪu�9�-{pe����MF߇I�+�Ԟ�裱�!g��"ă�EMى���3E�t��s��F�c��^�w�z�2'���1R�n^[�0}6�����(�����3]�.	4��H�4�����8m+N@3�>վk&k?�������CӒ�L4��OL �������K�4�������xւf�4�Ym���c��'��m��Y?*�*���yd����V.f��K���%h6��(��<�$�㖑[�u^b�be:v?"�x�(J�WL9�Ͽ��* �C(�n�obŪM/��B`A�ւ昹b��I��������a�%�A]dR��u�֏[Wݓ��/44�yF�B�5?i��Y�\J��?�T�"z]Y�;����W�13U�M:u���.7�oH]Bh�&~��l�UZt���:</Q/|�x���~�鞦�Ό H,���B������Ƿ�,�=U ����N"��H��ɸu1c��+���S��5�-�������������z�LZn�1�R�t�P�-�I�� ���F�-��#�or�h�\���[c��Ca�:�]/Zհ�SB��F����<@�|	���'�n� 2~y,�	B\X�z~ǈ��';�`�h�t�f����LB�����TR�D�2Ǳ4�~MWk�Ӌ]�{rw���x�Sϵvt,�>�,>��0��Z��0Μ:w�ɸ��a��X��`��s��4b�@ģ ��I��s�d�]v�\\��խAJ�6��;�Bse��K�w�U1��|�e���]:��pn�	S�ّ[ş�Z��;�E�z���.Ѩ T��=޶2��$�i�@�j�,��0��\x̸�f�X����³ww���9͢��B�������n�9���3�H0�E�"�:��R����w�+�7_@	Z5������<q �(��H���rV�'>�Qv�QX��%��ь�mK���Oo�Y[�V��"�,���
*������a�LfI}��P�.0K�JC_	`��"70s.��NB�
������\����N�a8�Ԝ	ʤDH뚳�d����P��{��a�.�Y�$�Σ�E�Rld�e|�}�O?�i�0ͬ8iXǷ�|���7�e�ĩ�S�C.3e˗a`%�բXw��v�w���I������S�c����m	�]��-�`�c�Gq�d!� ��|qI*)�zJHa!�r�F��9�o����w�:~��`�E�1�EX>;4��X
ڜ���o�qң�/+���z�&ObS�H�U��7��t8^�c����r�58JJ�M��Qg`���q�p�=��v�2=l�xN-��4M[��Ua✶C���;A��|����&B3��*���k_�HiҒ��'2����$J�J
H��E�dD/<����I�4�&@����� �HN}���IU�}�՛V/KއѴp�����Q�'�[�}>bX@`d9�_���X�!��u�������FM��k��z�_����8M�;|�w���BbyPI��i �(kO^�7�E�P󁦏�#�G!�7.��H7w4� Z�����N
�����}�Gs�>��� ��<��6����Y�x�SfU':���L�F֤?��v���Tm#z��̆�m��綏���"q�}c�@��}M3�� ���i��d��&�������	Ǌk\��VCF�� ��Fyɾ�~��7���e1d�<���� v�)�nk1��_{.O5�&�z�,T>
<�L�-G��!�������,���e��(h��m?y#�Qr�s-�d�^Z�e��fi�=�%)l�{�V��-D�w�E�Fk`u%���+຤JXD�b���M1�km,�[,�(.k��WW�HD�k�#��d�����޼�/;ŜW��A���V�:5��ѓ�k��ۗc���$,:���X��m�����	`�CB%u ����?��E�vI92E�Z��)��S��;��m���NR����,��2�x��v[3i2���-@�/2��i�����*�a_@!��;X���7:�J�9]�3��!5A���ߦrx����1�o��@σ)����ע�2���d_���TU;�b�Z%]�m-�Οi�5�w�ͩ=Zm&��a1�����毪�@m��]*Ru[9�s�5+'$bݣ�S��h����/p�&J� X��A�9h�T2�o�b땍�� W���YTA㵕.�Uz���*��	�st���c�).� :��"��6؂ʰ���7MQ$�#��v� ���_�,��˱住g
y$����a�A��uR��*��N�s �V��n�����)i�;� �ܛ�$s�D7��W�{�G]U�#��4ҰG}����r1Dp� �R��M�.x�̖���'�2��7
G"�nʁ�xq���(����6B :g%b&`~�j
8��J���@Ǿ���G�M�	q1�`vjTw��%߬��Tp��/�dg�܁O�M�+�n���Q����M��JcZh�rm�
* �Y@x-��-MBa/�A�4�Jb?]>ظ�4:���9`n���e�2�;E�ƽN���M���e^�j��Sa�::a�ɢ�:W?��2�F~I�Ӗe�tζ5�Dzn]���[&s�}E�=�`��MxP9 �Q�s�b"�5g�L2
Hf#�Y"�?r>c8�wet>�l+EN�d:�����>���/R�(Ӫ�����؍h½�q����FzՇ>K���~J	�r`RDk����S:� ���7HM��+�D�bs�4 <F�t��4<`��gW^�)\���q��:�>`G��]��<w�� '֕EոfJC����F�8�ŏ<�M �*�&��!1����I��i��g��'a�?&�2;Ϊ�����F�=�K���9�0wT��&�8!���k���VA^
gr�⟲缍c�^�"�9TpM�4s!�Ϟq-��O5U��w�c�"�f�H�<'S�K�:ym��ԃ��"���nH�
]�?n4����oh�{���:����5��Ԏ��$n�Dk�e��{�.x�	�}�{� �LU7��Jj���r�:FIۭ�h��u�'d΁O�$O��-��~������g�z5tt�]�_x�v�c�J�A�׏6�5��b�	5�o���4hg^:��F ��S ��z&:���y�׉Uh1��c�Pg����M"g�{z�7�u�G���|&jlt�3�5���FG��W���m�����H���盒���=��?d.�'Vyk�p`��7��o������^-.��F:~7��o�M9o�	/`���:�\3�$�3�T���*��� `�y]�O'��x�[�5�ga�B���7���x�I�D]�������\3u���P��Xdҙ��0k��e�.)� y"��(�R�G=�MSJ�Jo��:�NFFGضP��J/.��������-�6GYλ|s{�#�q�+����&������7/L���D6}��E�1g/B����K1�����f���8�X�鞮rp܌����+f8�d��t�Fg���w�kw�Sj�1�@\�Ď?������J��BV�*h�~ҰV\2���j���&N9I��N�(���^�⻿��a%E0���P����}Dހ��`����v��[58��xq�ǓڌB y�L�a\F�0IC{�W��0�vF��$��� �����g�ǈ�b�M�e�k���u=���Rԙ���u��d��[�lC+Ì��v��Sl�!HJTT���:N�zXB��@�єh��@p.U�	�PAuL�-K�7õ^'��/��.n��h[�Q��`��k
�����k���K|�`/��yn �3gA�yGw�=0��={֛�<؊;���ڗ]����sܲx!w}C���ݬPN܎�x��_�����gir(�a�g���a~���.����I�y�*�?�V��luďY/�H�1�w}|��GG��$���,=̯�8�J��ڝš3Am=�}֫��Pד�Jy�Z�拀���6��Iz��["���_��`��v��3�$B|s#�j�$O6�8r��L�������~j��&$Aw2�p���h_�R ����?�}%�ܙ�e�VDH���q���x	�{�t�vT	����:��䏐4��흋�[�#�.��xٜ������h���c'�����h��%۱غ�����c�o7�qV��Cϔ�r:�u9��Q�u�N�s��A���.�l�sG��^H���$�*�ExmH��ڥq%��V�$Z�m5V|[��Q1��8ǰCm��	cWР��ጻ<>|�4�{m���G�O�nWa|G )����*��	�+����n����9E���?��7�"O��>�Y�M\�Ĵ��:@ݢ���.�w�d;�>~	v:+]�龣`����ܱ±c*������]hB��ޑ�w ZK ���0,y�ފiQ{�r"%<��5�Ͼ���W$�2�#����(����<Z�1��C�6�ŭ��)׀C�Z�#��#��� ���rb��#D
���N�b�cfML�EX���n�J��車�o�'��! Χ1�RZ���; ���{�ΩÜ8�OHo$�ﻏ����q��N�������MBޖ�Ȝ	ԦN"�8&�sE!rs�1@�9���-�'�G!8mF5)P7�l������m��f2�XJ˛
��OK�[JTѦ2P���X!�C-������9y��$q�/Ef"�խ�Eya�eb�T��z|+�JJT��\�=�X�	�_1���$����� ���mw�1Q� �N��}�RQD�;?*-�g"��JD�jx� ���]�"�V��̵w���^��D������Q��㣙�V�q�����/q=��}
�l���#�*�G��ڇ�o�f �1����.�iw ����������Ix+	a��+�C�����T�?�3^%wd/�O����@��G�t��}�Hp��`��F�K�J~V��e��X�A���F�H�j�'�bT��}�q���(0�K�f�f���9�:h�q���N�d΁����Pf�9X��LI���?w� i�A�Rd��$ޠ `4$H�,��
qȢI�Ⱥ�x��6~м��|�Ê�Ep�@p]����d�-�~-��=��U[�Y}����)��9��o�h�ƭ�t���c]J�I����'L�yn��>$=�n����$K��sI!�6�h�U��h��������~W�_H��Q���0�v�9������Q��=��Iy9��d� �'�ġ����B�I	Q�a�pZ�pW:3XKɾ��������/.�Ⱥg�a�W�&1^CUS�hl�!'�i�"ֺ�tL8��uÔYV0͊��J����ؘ��|��+��P�H��g1a"�,��b�7�JN'�B�?��PD73��K��/���U�\���0����H�C�4I���i�!FfY����mm����Sx_�	ȷ� ���?�g�ˍd�B1�V�ôŏ	�J��9خ��I��Ni���Z�x�� 	4T��-/��۟�����ڋ�T�,��8A3V2��坧LЄ����t�P��s�{�u���UڣԌ���F�%(�	��8!��,qm�X�Ȋ"���p�Y�����bz��s<�>��-w;��Z,�!��>-m¶`m��N��}l3����E�(�᪘w2?(y^v���� �b�¬�e(�|�t,M�N{x�B�H,h��V0R#Q��h�4�YN�uD���(�5�<r�^5;�/2����Ή9�#�v���\��;���9�a�y�e�h�C�|]��mYM��$��FRoTT���ƒ�������x���У)����շm�A>������~�����*Fd��b��Z]��J ɟ��\�l��@C%=jd����1��h�t��8LD`L����V �S����VQK�[2�ON.��V�{)��=�'1���_�	�����b2ee�����.3�@]�k�i���fw0m1hK��ӭa �^��gj�@�k"���ֽ�������� �$5b�0��M�Z�(w@�pا4��D'�n{�b2��; f����qDz<|�eR� �h����sf�P/�{�a��dD�
Ua�vb�O���X�!�@
ދ����u��4V�fF3��CAIZ�M��������S������Fb嶏-#�5��GF���Hm�Ӕ\���[��M��-/���YE��-��:^2�U�aCv�L9P����J���@&�1Y'W࿙�AƳ�L:��w�|Vp��	Ɗ{�ܦ�V���?]��n���4t0���=�����j�fr֗�h��T��[%��X�T���'�4-�+w�z��uk.1n$w|9�8�8)��Oh����M��m�A|����z��ϰs��_��^";I.G���O#l��A��í��}%OLt.j~�`��ٳ]I��ijC��$�B�i�EMA�N]i.4��j����J�����D�nf���T�}��
���O|�ܡ�UY���V���7�F�/_½�:p�J��6A{����B�Rs25���E�C��;�w|��~���8#�9{e-�:��Z����;�m�_0�֏�`#�PhE��#U\-T��-(�G7'�c�@�&J�^kFGUGH���2H�qz�f�?��}��Y:�C��)��,`;��֚�����Ȯ]�b��B锩�;���Ny<r֭Bwÿ͜�M�M~�0��=byœ}&��ڕKރ�8���\��q��L�Ω&-R\|��d�D�H��뀷���ߓt:0ݕL�{L���Q����.f򤯱p�ۆ�b��)�)*�PV}u�^W���# ���H�G=Vq+mOAv_)O�K�F�P��7�$Ò���'��F��+����W≕�������Ĭ@I����'7�ҏq���0%'N��CV�$]"(p>�x♕Œ�f��^r�8\���v9�&��s�j����w.�G�/���Z�26hs�(��#ôm�4�y}��jM���R3Y����/�]�_e}�K��M�_����шك+e�͚B�O�����HKCET� ;�d2.u�o⧒vѪ����@�װ+m��]�:J��(kh���$�F��.<lCv�Q�ӖF#C�9''��lfe!��W�"�z��lc0 ł�t������
� �����4���r��)Z���1E�ң����C�.^^p{f?,B���3+�}��	ۦf��̆��!p�+��c��e����P��i:�쵒��^���Agj	�,���,С�Y�I�4�!G�V&%0�[9�<=:�,>t����¶p�qn�95�������� �C�ar��{��/����r��MTs�������<u����ޱ�i������:7��#P�t�&�*vΑ��@<X����������s*V*G�w� Qb҆�/��NZ4�ɷϳ_��BY屼)�C�O����9k��(7��+�1�Sձn|o������|���9A��S�L��Gs誷�6q)8���j�/_"n11��d`�Ν����I��i�Y�F��o5e�{m�h�y�|3s*؃�ZbSB| g佼$}� z����̋��4�;����D�C�����$G/�p�]��X�S��c#�[#��'����M�:�4#C4�M�\!ز3_�'�a�w�b��
J�����d���(%�E5)�����9�j�.��"�n��OVAS*$SBfᢻ��c�8�V]`	Y��`� .���-��ϕ��|�?c��h&Q�PPKl�Y$S��(��D�4�㎶M'��p�Yh��"�3ǜFDL�x'�5�H������������Y�Ln�I�T��&zm���1�����~N�=D��?d�W���}���4~��z֮�;��R�M(O'W���d:�l�c�~L�mE/6"��a��ؕj���4�a�F�����A�;� \�ֳ��R?eL���+�X��K�����s����x�G��5@g�"�H��}�A}e/��� �RhɆ{�A-'�K?=�l�&���ꖵA�~��z��J>\�U@��XZ��,�'�Cʑ��C�@�f�l���;�g�v|����f�ފ���|(�m�����C�����|J�"aյUY����^j�+?y^����!:�ģbRi�B�ޫ~V��z��{���׈e��x��0��N�����q!��^Ĵ�p�y�3c���z���%@+j�q�r��O%)<eu4�?��ȸ�XGDi��[7b�Cg�ŕafC7^��]=g߲��:�BJ/ ��'���J4`�C��Հ�����d(�v̸���C [�7F�L
n�� �f����u�QV�%#�8�����>`og?(�3�����>��p|~�|^�$�R�y-�e#��b'ck4Vi�Z��{�;Nv��5��d̆c�gR/��XRq�!C�6"��"���KL���v�:67J�����A8U�sSw�n	S���c<��34�
3j	jd~�Č:��l_����θ*�xy��r��^6i�A��������-��U��3	O�{��t1Nc���n��݊~��A�S����� ���/RM�p�k<��~���P@Z��NK_`�@��*K��* ��A$��.xG�@t��d9|�>/��a�#_g�z��Ls�fZE�n�2�BHMz��.�w�]��Í+#��\R��i�f��pY��e�.��KCپF�3��(�ƞ�_qj�ҩ�sCW�v�kZ̤����(`�$S��1���D��J<�k2wLr�EU(��ڭ� ^v=��ҕ>�+�TdTɫP��o��������� M��M꜅��M�=Z����}�_�l�I�����[�������r^��n�&:�Ҙ�:��PIqI����������Ie�܂nǴ�b&�/(���Φ�q�ĎI����~@Y��`�{ �`���E�1N7]��*v|�Qd��PmVM� lԱ�j�R�r�LT�@��~�Q���J\M�K��ۨ��+���:�͋��(ݒ�w5P�0]�|7`=�t<�ڳ�9E�P�����߄��û�r.���PO���l�ӑA�+�O`6�4"�������tn���[��\���Y�U�t ���Y�d�����R��y}$T7�E���>J{�a&��:�l�����v�j�K�SP���"K+=�A̋<��7>i�5�H���܇��hq|-N�w|�Iit�%�K0I�Y��7�=�s���"��l�2#Eu'�F��A�.C^�WN����+���E�χ8��	/0t�4S>�@%g�vفG�w�2�N����L\��<�aG��GHh'�	���w�_�����-��i��-J�������Z}*���|R�j����eܧ���F<�+���MB��H��(mXE�;.�|O� E-}Z$�Ï`�(<3�g�+p�����Z�U�	E�x�h�-B�STc:��ݏ��dZۄ1k�Mɻ��!ef_�K�/(�m?�0���}�oeZ��cz!���=��Zu7��|,M��9L"+�#G�K�eH���k���8�[ ;4��h�;)[�F�_�p���(#E�0�7���7�UЧz����1}����I�mCp���и��r��0�(Zݦ�����R;�C��X�N���B2*����ǧ[�X�:ƞ�!z�P;U O�U��.�2L��(�6�C�o��o�d�t��������ճ��X> �T�U�%�F��p�@f�
৤7 ��a<��Ԯ2@���$�7:gb�)�C���WF������gx�W�N���DK$���mG��v�BH_D���8�=8+�T�����[CJW����V���*uĒ��MD;�t��+�(����E��L*v[+H�`w�x#�P<���N+@ʝxŘI%��k(r4�? �-\�:�e�*C*��W��6����~�m��f|����Ayv���8��[ڱ�V\i��M�D�08�s�~��%P��/�.h�c )�"9�h���H�A[5����H0�Ҝ��B��7.�(�"
���;\�¬����XlxV64EB     733     250ڜ�ڒ�nL�K\R[����m��KAV|��V��a8�7<�qNu�eB��7�����h%�$m@p�� �(�X�=���ˢ���f���扯�p��q�<�V/�056��~&��D�u��\��l*2�c���V�p���6�n9r�`��k'~Ձ�_K������u���P�T�Aźq��(Z�_�.���(����[�O����]��l�6�H�k��~��� ��<q��Xx�_�ï~Y*,cl�ĭ��Ѐ�sWo�Ժ�0J:�("O��Ԯ6愿� 1+��v��|�9�|�~�&�{�G���CjD/�e�Tlw� $�����!@G�&�7R���kW>crP4=���N�ӧv�Č�v�5%<���wX��Z�t�#�r�"8i|E)�4cG�%���<(
����=ʷ%:��A"th�2�����:y��-s�������s:�7\ �	���#��WdE!��\�I�G�|�(�&���;�_ڦ��{7I:BF 1<KBŹ�b|4S�٢��[!]FS&@��E�o_Ney��k%yC�nduU}YW���(uJ��X�������>*��&��=