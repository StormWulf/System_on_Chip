XlxV64EB    4961    1410��(���C˗�ř�Pb�S����7X:ܔ��6�.��xNI�=A.�I��ѥ�ٳ��h���A��NvQ5q�b�0C�W|5��|*�ӟ�95b��*�s���.Y*3m�^+����O$�7��?�X�0t��p7R"�'	�6�a]K��Ae˄/�$�xs����{���Y[?d��1�G�_m�}��2o�=���b�D,]���R����zc�*w~B��(G-�~�%�U��8Sߣ�A�di8v�.��_l~��7v�
&�H�T������$?��|��)j�;�i�n<JT*��at}z���C��IoI�Zq�*����!G?dFS$_���]�]�s(���Q��۱czR���Z).ve��� �=2����֓ʹ޿������<'+�H%���f6d�Eh
�z�
j�ī�"�h���	d��?������̢"^��<S �%��q�����iyk��4o/4���(�R*�]��B�R��2A�Y�5{��A�c.A�	<̱��Ӧ���^i�!��B�"�΃�a/��F������ST���% ���ZN����*E�h�����7fЃ�8�!'٣ �����!=�Bha���}�~bi���0�I��q��}�Q�YN}�v1;�V��RR��i������=��&o��[�B�����b/�Ow-��\�r�z��{g*A�G�mcz�h�#�侾��
4�\'�Ζ�-�$������}�wĐ�(>�0�>Ƀd�<�Cjl';��r9*,B���9�Nc��%��	XE_JV����Zx��~���z�qW��耹�kG|y�A��hb��Crm9W@��d��"�v}��8�9���ŉK�J�@�D�7ruF"������u ���1Q(P��[�N���1��KQS"jոn?��$�uI�Dxs�`3k��y��Y�hě���������G��m�����M����*� s�Of�];��+ �J��n�P��A98��U��H�y�nC����!�u��Mv5�î�ǯ�A3�}:�e�+���K5U�����,�1!�1�8?���;�>���tO�7y���
6��dSdU!;k纑0d��<+2�����(�����L�S<����m-�2cH�x��S�^�zUE0t's�,<:��+�<�z�c�&�t(nx��2��c�R��u%�~����B[w�iH�\���l_̳c��	U����c�Ξ�&a2�'3�D�
N֏":�vC �U8/�b6�/�L�j��H��Ӻ|������Xk��%�%� �_����`��޼2�%z�C�e��;���	��V$[�t���%��\L����K��8t5zҳ�7r!oK*O{�%�jr�S��������Gf0!��П�����s׉�D�.�":���{/B	�����T�1W�&���Q�S}������]���5K����X%�t:H����1���3>W,���#���4��4�=�|OFφ}�aDG�>�e��t�����t͐S@�R<��;*��-G�3�{'i'�s�k=����+f������+ț�'2�kvJ$~Cwށ�K��Wt��o:hˢy��\�8o30������D��F�Qk��	�߭ܝ�w�����G:r��nk�B��3IO=�t!p�,kFߔ��wmq�jzfs�Ȃ����/jx|[�7�Γ8�XMB~�?J���ˎ�=��<�I�[dX�����tb=�Q�#�n��\Z�Օ(3|�DQ���$���5R�<}k��cq�l���}�kjz-�>�H�eJ��Ɉ�|	��屇����܃�����	#T�[����$C
"��NH���c�dggI�v�:��-��H9����bu��-���J3�����:�#/`����F7�����uG��`V� �0g��)�~�LXn�Ӻ1�ƞ�1�Y2 �zCc���qB=��b3�U�הj��-����4�UY��a��~��6��m�5ς&a�ܬ�Y2��P�v,�AD?���h�qy4�as]쓺�������.ނ3��	��#�P����2�8O���L��Խ�R
���GvYI˱�#��nAR��P���P�^�G ��D�/�iL�ú�=�+\����7��hd�w�]8F�Z/H����V���xT�����t�0��T�'GRk9���<t6IPM�)�.u�̹��[z���%�7���E����B2�f��h�� �BF1�j=��Vu����eO���cGc�o��_]�R;�Ƚ�D�'�����i%^�Z��s�)8b����\X�\)��`5nq.z�:�H�(OQ�2��h�o��p�d�����X��I��O֕*���C�lzR#����������U���J{j�nܸ�4�A�c]��]��ُ��nH婂�Mҽ��aF�Lhq��F��|�)�2J��_���g��&��Q�����:>�U�mb��*p_<v
�m�'i�E����-�=�-."�LO�~�q�Kܞ�R��2��S�ɗ�H��;�E4�x�,��ø �B{N�BnsDNkF9�B�C������H��a<S���r��D@���$+�{�<�POg�Nbg�s ���˷K�,考���A�9ꖦ7t�S͑@�ُ��׊$�-Iޥp�0/��vE�I#Pp[�ꈕ��%�-灕��`��t(�w7r��ZȈP��m�c\�����^��V2���%��
�$��D*3�H�T��e�uH��re�r�Qg� ��f�X�Ǌ�7��K��U��X��0�eM��$�gmR�	��,eP1)�%ו̀hW�'��Nt�ՎN����jwV�~=��.���<�L���x�ѽ?�:�����h����Cj�e�F$��Ii�4�+C�'���P�|���G���l�d��.G��ɽ}A�i�G�o�*�.B��Sp:�g��T����� 0<m~I����6�_��0-�ԛ�~���1_5�f�M�����N�nN�E3�-��%�L�*�T7-���Ւ���a]��F���
�Xȭ�M_�G��8�ڈ&{R�0�qkT�e�Ѥ�� 9� {\�pq�He&&��X^'�ؗ�vT�9XU\1���9�cJ|�k�DZ("�+�^=����"YIQ)�
	��N0��L���^�ym$�+�ψ�Q#y[y�i�N���=�(]�lS�HX�o�o����o�,B�+K�I�Z�����D�ˮ�$���N��h�
zM�Ҕ1�aQG�n񱕞+�{�ߔ-��B������E��)}�Z��������	�����鰬<H���&�$o(����C�`�y�[:�u���;���S�#�V��j�6�x?��%��8s�� ��@�lWK@���+}i�/{@Nl�=D��HX1o:}��N��Y�l��t�0� �y�]꒤�m2�t}����U��ƫ*��a��@���$����t��V�eN�Z�-0���t��0��}C��2 �܇�^ ~{�4cֱ�C���at�����e�@�A��:����:A���
�M
DE���
·�-i[���Tk=R_��lݚ(k��`��g���D��p}�I�N&�yF��Ǽ���y6�15K|C����6��9J"i��)�
����m�-
�Un� _鋕
%��aq}ŀ��}���Tj?��N�)�_�~g�M}H7���]o���hݕp]H�F�9-��%nh��˲]A�X���Sc�C����J=#����-k���Ű
�b�Р��Ssb� ,C������j�,����믊+��[{x�j��	������$DcS2���̛嵐�p�0�"��~���V��Ō��O	V������ȇ:�����C���˦��O�ۥ��n�"��:[?x^���k ��+���!9������� fK���A��Ұ���ay8�D^�zB[	n�?|��s�K���8�o�eS+j�,
�TȎ-�$�J+7�`_aAt��͘9|cz��t��&c�h�-_"��^m��4��^�$���@�֯M0�O�O�Ğ�[���p��  L�Z@����KI����1ʺ�xWvI�$��,iP��ʷ|2���� ���]p���xU��w��Y]�fE�f�$�g���՚�H%��m��CJV��ſ�ē!y%@&�ؒ?����(ɉ-Y}_YxK�ŗ11��e�� ����y|w^��t�ݧ]9������@Ŕ�9ө��Ejs#"Ѝm�-�e@5-�~̀�p~���ӂ��Y@��q��z��#uzG���Y�;9lmj�4����IˁB�>�n�D 5]+|���� {c=�hT�t�n[q0T�Ym��(���)�@YBxη���ģy.�Yl7�hR�v�(�Q(�&36�߂����)���He���p��׫���q����,�o�y�m���"�xML�5o(=i��5Dh�
���� ��lef��Ȝ�A�E��i�o3T0����@.D�޶��ݤQ��h��V^|�=��[dɊbo0��fQ��5��)mkb�	U6L�4	e�#�������s0�i��6�y��O���L���>��^�It�.ֹ�	3o��
{���wz�ب�3��k�{9�R%��8��i�OE	�Yb����@_a6u�_F:U���S����QmD�����6�jB��"�C��J����
l��_xן|� ��W�V��J2g�j����!	�@o$�-�����q�q�[��"�[�l��̪߰c7��KMx���Y<Pɶ�>ڃǠ�c���Ͽ��sP.h"��+%�}��_I�J4Fō�t��	:��*l�ZD���J����e�� �VhU���*ţ2���䜑� Ng���+4�\}�������/��>O�L"�����Ӗ��˭,���{�w��ҭPA=��DH��6�I��}�+ܣ��RRfNŝY�JE���5���-L�أ�������J>-p��u��á����T���H��������n3b$ \sidf4�Â����ȸ��9�媡�F�?�\��P���:E+�{��H�	epL+z28�uvYq���b��g�