XlxV64EB    1e37     a80�l�\�J���@21������	���~*je�`����n�뱉�]�˹�`wb
݉��$Ԣi-������d/�nd��9��S�4;!�|���cj| ?����s�96XeYx��a���f�������������]��)b�D�P����./x޻@�w9;���0.�-c�c�6�4��WVbE	���m� �}q2_wܐ{�/BEV�-d��Ro�S���)'�>o?�5e��5-�G�;s(n�K(�6$�K�Թ;@��)n�({�������Y"�r�ˮ.�w��Y �f�� ��?���-�=>!�L-��}ܟ�����k���k�Dמ��ۊ�.t�7������j� z[c)��	/1��Z�_ 0s�+��ʽ�����wɁ<2������\��9s������U/�pH:u�!M�ۈ��-�4�t["�{��]={7'�fE8F��R�*�)G.�&�<w�A����j��i�IX7�lz��N��u8���*�G�H�/�Վ���)�t&3�b�'�7���ϕ;=& �T���$" �U�{*>�تC�����jFD���]������ͤ����|}D�ސY{���?�qv����e��P��F5oٛ����t��Hn��t��% AL�Q>	�z:�J�4^:�c�j�"��顃.��\���&㺻f��D�#z�./�^1y��G�ph���#����:$��,�.�ie�l�T���A��
�����a�
�Znz��iSJPtI��� �C�q�Q��O��JD!�HD�d$8��܆���� �!�yj!X���M�@�~��|wg��2�����WːR)�*���,ݱM�9�$�g�Qr���nf��E}W3`�w��t�|���h�%����Z~�ܹ�@"��=e �N���~�ݴVD  Ǖi�?���,à���ET���lς�5��)�T�x�{�uk��i���N�>�q�υ�/)n*i�nzy�;*R:�$�*H�(����@��=�RAETOa%W,��!0���R��XF"�.�c���2*�j�+w�$�Eك���T/?�%�qN��,�����e�%�����r+)J�TF�1W����6���v���`�����{�s�R�P�[Ǖl�\.�5��`[�H1�� %c�^�ލ�/�ng����X7F��D�.;�7h���7U��Mõ�'�+g��y��w���CP�g����%zXk	TXj�����1�X]����G���6�����SSJĻ�|���o���)7�r7���I��bVd�<���n'"�[S��"h���ز;~Z���^�H����ϳ��P�����V.u�RwOւ��h�/�N�q�x8P��0)U��ۧ���c\ɦ׆>�Wa�h|�<�j�<䗬�	���j?؏�a�~a���&rЯ�("�DՕ6"�I�(ikC��0j��)�Soy��WȚ&��Ťh#wi�3>h�т(a:M� c�޵Z����RX#�w�L����Hٲ$ ��V{ؤiVsg�)�/n��ʲ�!�6�2Ӗ���N7��� ��M8{M���.�L)�/T�-�������%7��n؃�Uoq�̮�1��ၼɥ%�>]��y�0���z�,�B��C&�v}��2`�����/�"�M,�zrk!�z/�^���+�=�xq-;�M�$���� rÚ��T�]�S�T���5a�� _�◺4g��#�d�z�tmK
HX�9�hV�@�=A���$q��j�&�����_��27�-m��~��g֣u @��n8SD N�2�8@*>�i�+KQh�d�l�)e@����D�S_;�oP�u��3͊�� �H�t_R���!Zr������B�V����5���14�/�AU(��H��_V@7�'����N�YK1]mP���i��گ/Cy�6|'o�4Z�|�fwt!�b����]}��.e.�r`.|Or�16�Oa��)Z{�������V<�GX ��� ���}�	r�%�:�u`��=~+��趗YQ�(ٞI1�6�չQ��Yzκ5��3�\Т���q��y�xK��#���"3@=��cg��nG���Ӷ�^0�����M�����j�"X��q̭����	�]���@���[=��)(ĝR�~�{;d�R�2r^���n��L 0X��#p�S{���8o?�0��!��G�(��^S4��~Ф��p:�|�L6�|����L���g�{T?�L`"��G���h(�/P��tַ��bM�}�!n�o��@׎7��� ��'}�.�tS����c������X<��|��"�$��Z]��h0od/��{r�@o#��őϱ>(J=��zCM
�*/
�M��ɿ`����MQ{�"�Y+AT�*���ӑ�p)�ᒄVQU	'�ԝ$;ڜp�Y\�ie"����������Z��m'&�yq���4I\[Ď�]46푄N��'Qv�_)�u��nc���4�sS�����u�8����Z�d��H9�1U�Y
���������A"	��>��T:'U�B <����c�94�¯�m�`\x������_}��������Z<��}9�6A��3���-$���Ԁ�������zIwD�1� 4g ��