XlxV64EB    3f83    10f0��,���"Ը1y���p��-t��~�p�;8�b����F���Z��v+���f�4ڳ d�0c+�W�U�!���[5Z��eG�GtTRk�mo�b�NgM�_������9�}��ީ��z<R��wF]��eWP�o��j��Z��	�=`���E7�8j�Į�f�����	��фu�i��BD�U�3ɷ��7��5;�U���|�$/X�;�p�x�=[��뙙����b��� �M2�J������ù,�� Y�#@AiŽ�y���J���td�����|+LO-�_?:�Pd���W@��x�o�n��7�$�Sh7SЉ��N���D@���)3�Pp�%��<�S`��eM��\���28�eIO�� 3���.�H��ͷ���Q������1݂6�"�7o��_ԛs�-dk�b�r��ȁ�m�Q��k��	�'�s��t�+�8l�ڋʩ92����4�
�A�����2PB{���Ҋ��]ӂp�SI$���.A�_+��O:ͩg�m�;�[͏J����Yh7�g-/e 'y�9[*��ß��$.C�$7�K%�<Un�+F�� �?6���W!���O[!��o��f=��?Ju�G�T�
��T�s�6�����Rb0d0�P �#�����ow&\ܹ�xO�	%脜۽����������nƌp�Q���Kک|'lˋ�o��C1+ Z��j��^AuP��ѡ��v�Z),и�ݡ$�0�����T6�?�'%s06���o�~u_?2�y� =U���LXlīR�$��Ș���G*]h�fa#`��w�6�O@:Rg�7�	�H.`0�HC�Ǐ�m,*��կg_Ow�fH�d�sC�������`�v����t�� �@F���_��Dn����E���T�6���ﳡD�Pu�wA��$�����ýL���"}�Xv�I
W4���
;�4r�"�>���_{\��a�O����Q]���?�ys�'�y�8`3�a�Kp|1��3Tg}�Xsr��G�H�-O'�:9i7�1����c�I��!aF��qФJ�V�?��"���o5-Q`ú��[�����9=�[O�D��j�ȌҌy�����X��<���u\�ULH��	������X�juI!�%Z�����a�H~-��
2M%���I1?�����jyيm��P����q�-_gm_�I�S����ɛ��{��ci��5^����
��]��1��ދ���k�C�^�u���޵��F��N�f�>9�'$�����r���w�l=<z�_��.B-87�%�lݴ�^����&}��r�/B�?����/SUvFɰ����MK�g5�y�'T?	�������Q��}�?]Lv���Z�Q��Z�Y=��H�3�V��:��v�X��ڂ'�Ý�+8P����K���­�b���j�20�fU�Hh��BK�D�k#�C�U�kԮ���AQ��c��O��1g�c�9�v=Ó�L[S�pb�i8N;6��^C\V�us�@~~I�^/�����ݽ>/w�ʖ���;)�d��^��k0�"����"�&���`)�l��#T�}����ɘNj��߼�C	�a�x!�	����܊>[��և��OC�ٹM�y��{k�2�TdKz���-�6�N��*so�w�$��vX91���#��T��4o�Ui�]�����ۥ�b^(����p�쿴v\����췗ag"���uU2B���=��ם�\;b-�	'�6FT86@���hK�Yb�^�rP)#� eg1;��f``�%d=�g�)N����Җt*(AET��T ����;� �H+��B~�J[l�6���I���R��T+���i�5(�E�`&,j�5?�O0uƮ�pk�c��!��$���)�;0A��]������v�l�O�{�)#;NH�f�!��QSv �&�n��xx����<{���Hu�])؀�&AYW���QwI!E됅����a ^�e�.W��O�l��`0��2c���X��q���ɶ���۷�sJ�ol�T/Q�ꊃ�J�uf��TCi~�&P��l-��$����#����aGpa�z]U1\.v��A��L�x
���&��ݶ��V��T��q��36L��L�!d�T7�>�������H���g��;�Y���B�l�H�̞EA_��Y&����@�Ԏ���&�#H��l�v��g�f�u��t~w�^eⱓ�D@��Ub1�F�d��=����1�E��Z�=o�~�3�N��o�.\A���D�:�m_��I0��X�����,��s�b-8O�`"l�D�k��u��=V,Q�K(_��g8grDUƌ�([�����C�Vy��f_�6��U�ޑ�3��0o�D���L�R�E���Q
��t�`��bq�ɝ���|����S�*�;�$��,��f\�+�oe�=��ٲ�f�D��jtI�퇄���|��[��O*?�u��l�"?�ħ�� �.�����b��R��l��ߚV=��FbQ�x������ ��i+d��JPsa��#�Q9��b�r#�~s�/(�N#�M����di���^��]�g����2̙�^��2d��B��^��ʟ[�0�M]�uҮ����p��D2�U��j�AEQBDǃ_(��p��Zrx�,NO �֔Z/|8�6�b@<������@Y'�H�1)�S�[H##�܈CT<�$�2��if�w�5���[�@O��K�8��������D-5og�8@�t��1ؾeʝ����g�u�v'{��n�����8�e�
�Vh��i�5Ѵ��3���۞k8�w�H%�V��|�M/�0`]�l��w�a`r� -Q�	U�}�\8렅���c���(�Y��� h�� ha7�,m�LU!� �~��XӴ>i�rW<�ND�����倃z�yi���.��f�� ��@F�M��%��ҝ�NDS�J��>{#?���v8��w'`>q�^��I ���lv�n�Q$fŅ�38}�KΈ�[LMե2�Q~��o�^�8<DmB������Y"/�LKa��$���b(�K�|�5�|�� 0>�E�,6�V�C�.
k��M��_�jx����N*����q�62Wu~_H+�R�oʛ��@�,��4�q9>x���tR��&R@n���F�9�(!5��?K{��2:�Cy���h�=�^�Q���[�C�9���ò���@�ٔ�z�n.%P�T�MuYP.Ϯvg��~���31��?kT�޲�x��~ ���I��R�.�2sd:�̼Vv��U�=��V7�ˀJ`��������<�1����ݱ�Jsi��r���])�{h/�ؠOƾ\���,��z�`}}�d�:� �f���?��<tv'r!��^�&he�K��<���[��Ԟ�d4��=���FL�Yhf�ļ`���Թy��<���HUsJs�GT�>�w�~�א����R��a�lꁫ�ۯg�[{���?J�·�2�vw�7R��^���P6%9�r� ���0�0����%/�$���Y���	�ec!����#��A�?�5�T�/3w-�l�O�58.DI
�!��|E��;�3�*^G��7��bn��]\(cY��������A�J�F؟��`�PN-��d��oi�7���/{������o����q*�7��A1_C�a��;�Nz�$Ӽ���rEЅ�0��o`TZnD�7�2B���v��d��ز��*��@Q�P$tP�w��r��+��6�+����>h��Hk��9�"�$��s��H�t�yK��Wymp�=̮�����eߝ��H�>���?�>��_��x���J����Û��Q�MT�2_�=.�F䛴W(H����\��LnF&,��/�����g]v����3������)Ā�G_�"j��+`/A�gޛ���Nt���ܸ��_�q�y;pq�� ƵM*��%��{-T��V]���ؒ�@�1���./e�hG �8�%!0�L��"�d���g�"�i�9ڦ�A���O$,}@mXs6���p,L�~��Ԍ�X�_�w��1�L{����&9{�=>/v)/��z,p�����wHQ,F�6f�+����̀:<(!`�X.�)�^=�9�2�x�7�zN{�`G��\L�j��Z�A����^���#�䀔<�r`���C���S�LFU��vI�<	�wZn ��r�����/F��(��m*AO���%Źؗ�u�{�OB�N<�H��QXB�V?Z�=�2�6&���.���&o+}�dS-c��D6��9T)#�E