XlxV64EB    88a9    1bf0����{S����/���mraO�cՍ���� �@yK�0�9rF�L�1Ϻ;3n��T]kŋ5a�Ձ�y�"����hF�Ƀ�aZi�@5�W�����2ye0��t)$���';��6�ع�����}P��ʊ�Tp`�����輊�P��xU#�!��&��y�����3�{JSdN�L�0�0��c6���n���q��J�
�;���y�I$g�����q���#�y��)@��_��߼��c�������K>��,ۺ�����
����8A����	�i��������"V�E�me\��/=�kT(���6`�����^d(\v��Q�p��a�b`r.���^"&�"��2�)����ޖ�/8�u�3�eC���U�7�3U�G7Gys���Dn6ӎ,s�����������K�]����=����T��$kɂ]L-��"�4S��̤�`|��Yy��ad���n���1+xè|n���z�o�sT&� ���p�o�s �A ��#��27Mp��%w���ga
�ϕ����4Y�Z�C2e].���A$@vF뺑ٓ��V�}��_��R!�����k��:��67���'jά���?��8�+�|[*ÿ�DHD�b��+<���-� �~r �
eN�va�J�5Ky��Bތ�1���t���`4�C]�e�n�n
(;>v���*�4�$E_*Z���Ѭ��Y[;ol�Hj��/o��A�]�j�n��	0�-�����Nu�!' ��"�4�!-���hX껕4�-�P���8H��l��)�j5�L�x����A̓=��������=6� �!��u�usp$��"|���Ӗ�͓uF�wX^7RZf[�Ĥ�~mV�K�K�U�J3��E59`�B��E]]���sʢ�6��7�w���<I
A�cGa6��Z���-*W�3�,I���UEv�q�@sdZ�!��7�(�[��{���4����<��(|AtA^FC �r^��{Ⱦt��!D�(;�_qcm���t<⁹��[�������������X*�	�\��K$	�
B���T����|����I��R���쬘}F�zx����[㶨�D�Y'F�ٺ!����Z4\<pO�w)7�b����Q����-iЭv�p*�=�ȿ�\ʣ.�~��&�Ѕ���A�l��M���BO��1D��z��vp1�=G󵏐�e��$�W����Jy�7�B�6��J*I�f�3 �ݫr1�� 3t����,��y�����;��B��[���!�o�r�'���9�~�=��j��5 )n�#/�/���@����凾� ��g�����T&�.���E��' �XE˾��U8���k-�
H�F3f@s��@�x�����.I����4u *J�؀O�'��_S�I��tD
���X���Xv?%�Ö����
I��ĘZ\��������}_���K�Ch%��C���,�Mc���.�{�܄B�L�,��a��b�2��a�Q�X�g�J�8���x/��S����P��<�A����o��_��>P��fk��+�U�3+��`��5���MG[�:�?���o�SE���?��S���iه�l8�q��1�l/X����k�4DG��3X8�`��@��T���J����U�R�X���}��ߜ��Zt�P+�@)t �>��vL�H�y�diw���ˁ�<�Ma6
K�T(��EU |JAR}F'?�`�h��mtT�\y�s_����ζe�IN��EzNߑ�f�e#�,<�k_�kR�?���:�Z��l��Mj,�w&�%ƈi�I'@��-a����u���� ��e�h)�v��1�4�\4��T)x�J�Gh�y/�(]�#����?>�)�(�J�jm��R����l��1�����0�o�E�D��kv4�?�ci|o�d��{5��;-���.hKK8��L��%��I�����Q�ҳl��t��E�S����d��z��y��$���'���>���T�i�a�Z���֫R탍�׹}o���Mv��|��w�:����F$OIN��[�Nq	���d.����Z��Ly�w$�ӂ�����B�Mtp�6�ED{3@�ߖ^ �/mB��K	bF�^"d%���cښ�]������m�h���࣑�v��;)Y9�B�KS:��'�XHĵՀ9B�������R�Ή;1	��ms y�[�繗�s� � ���t�i���sȤ�"�T1�2"��2�\����5dj
-�b�[�og�*c��c�>l�cnp����yn���7Q/�<�[�=Ձ�q+��r������]y�9j�X�,dn��W��cH9��m��ޥ��V����*ş��N��0�����&�#|���P��U1k�׹�h6��h�쪆L@��v�M��7h��F���(�I��l��ڞN��J�C67k�ʾ��Q��%SP��Ɣ������x��b��&��>_��59�/5ҋ�	��H�)�F��$��&N�rT���+�!z�%i����5x3�#m?�K�6�(�,)^��2e@YM��7�������Ӑ.�TL�ס�)�
��Vv�CyD����BdEp8?�\�o�ޫ��~�?=m���`��tx�y�G�s�1��ߒ�v�>q~�4v��Wj���b��X�Z�|t�Om��>W[���r�_�g�r�_����O%�a,�#�e�*�e;�5%����f��t���|E���T�)�d|���~R�2ʨ 8L5�!9
�����]`�'T����G�&�C	uwEy.\C��>Ϧ���p�Sػ�^���j6�&��Wn7�E��c7z�t.t�WS����h
���Je��A�I 8F^?��~����N��oq�߾{��6��B�C�?[Pl�`�AC8�-A7�	�T0���ీ�$�9���|p-@4��{���R!��4�>��1���9~�]{Hu�� �V�����>�nXN~^2���A�eY7���d�����L`X|�7qw�/�}gҭ�����s�L�"�����&R��X�-���� �\~ǫ��9<�|Q��(��^.���͠��_�ھ��Ԧ��mTcsH�w�?�ދ���7d��>ڊ��9_e)�E)}v�H�NB�T�;��L�����e
q�ܪF�F.ax�Y.I{v-_�뜐{�y��40����_�ɦㄾ�U&��-_���ù�ӎTI�<��� �S�O�ӤRaphd���e>@	��Y�c/�R���3z�6R+��5�1Bi4Q4W��$�w����kK�>�,핮UH\!����
���I���W�˂�-4�ACS`��Jk�v` �8AO�%���?�D�)l+0��E}��ӡ����_���-؀�,������ߞ��}�� ��0%�?�D�{���W#5}[(��w�e�S��dl� $�(�<�!�^먩c�3�ʏ�~):X�����(aw�p��C7,�0���q��uㄠ�w�Š����|���mA*�������5�'���Q��C=��A�3?_%/saM�~�hp���zׄ'k��Tu�r��h
�K|�!���"K�7# ׭VDo�|K,u?4���`�x|��4�#E��_"�S/�oz��h�'�~a߀�m���s��%����&����p��s�MZhYM514a�s�qU���J �6�Cד�	��Ђ�Rl�yVh�q�������=���}L�2HНҴE�����e�_T�Q�`������Y�5Ys�x����J��M��ׄ"_4�g�ȃK�ґa��GQ =�x�fZ��:6n�nr&�K��E��"��0�戀o$'�����6�G�3�Ra�[����*t�UW�_�v1}5i}A�Qg��RRЫ��<=@9ߋ��{�@�7�7��%�2j5�CX�ה: ip��g���O{f\�k)Ñ�a�������Cx^��L�3��e�h�Ҕ��n�� .���0MK��#�d��t1�HQ0l! >A�&��F~ڙ���d�S��X$S.�&��Y��#5yԈ��(?V1R��ƀ9P��jߐ��8~�Z����[}ݒ�j����T�}l����i(�� �������E��a���=�	#<��3Y���0^�[ӳ�&e�������"����"��G�\��c�K���#�8۴�a� �><�E�X(N
����,y��9����h�������uC����۳۽�b}�YR�P~5� �ܵ�r`,S��8�N3��J>�+'�f&���'��=6��ե
�lM��o�U���)_�bN���0�D�G��.\�M��:`�S������A��T*���"�t�� vJe�3��)T�φKy�� ��XW6��`zZ�YЀ�x&����$�o񲬝p���h�_#�gP�ϟNLJ�v�� �ky|��416�]~�Q&Z�$) HB~���kө}2��4F�g#��3�Q�s������Ц�d��.����� ��l����k�H�F�S4tr�Cރ˫�. o|�z��Y��0����B�7��L��S��	�U�d�]7����:��U4�_����^�TG|Y֠l�	���IY�ٺ��&F�ߌC����XB�C@H����h.^^����Q����1;���$����g)��vph?�S2�&��(,=�ں�W�KTR��I�[q����!$Ki� �{�S�شk91��]�/#�M�TƾҖgd��j�ɼ[��{��!���=4�Yt���c����,�]Ç�A���-`s���%e�ΫS��6������=� �e���[j�����ƶ�a����%)Nh�5߿3��Wi������b?B�c۾�}c�� Z_�1�fIjn�8��;�E�9�8j�ӥ�I���Z�/�W�
�V3�9C�{���iV�q����J@�����<F}����y՞ZѴ�(�b/��ec%�M�r��F^��۠*�>�kbI � �����r���Y���d3G�E�֩��Z��H�bOr�����u޳��#��zERGʛkJ�;E�'�c	�8[u��~1m�`0�jY�k[�~������a��eFQ4[��R�Ln�UӃ�R���Bݪ=�#ۘ�Ո�^��K����>��}?��9�#�ϼiQo�=��_CE��Y1���n�Ȃ���Ֆr!�Do�,���C�Twڰ��x�n��@}�,�kDT7�Z? z��2Ѭ���+��k�A95�==)�8N*Q��qFT��Q���p(�"U�x!{�)�}�yB�>1n��\eq ��]1h8�h�BR/��v:T?,�/�X%�',j�T����d/��+M��+Mv���u�br�l{� 0D��GV�xPC؋�hi�J����a�U�iBf�� ���nZ�63M���o75ϲ�5fb�� �F�a�d�����m|�1{���P�*)�S��˞��t�$5y�d;nT�#��' ��|VѦ.�͋�Ɵ�yv
{}v�y�����,ߧQ�<�qHu#��ߖO�aE�=?�	m:2��/^���>R�_JARVt>p�Qv�Pc�<n�@ȓ�������Ki�	?�r]w��AA"����������7�!�ȿ��,������k6~F��� >�i��6��f�`�ӒSh�����/9Z�r�M��]�N�=H�{`���rEW6v<��V�Y9��B��|"��	�xR�:|�(C�7�P�N�`���_��(_�z��e�z�`��������5�������*�	�8����J��A�
��#&o�.�3 Kc��~k(�}r�C�	��k�����8��'$��e����vv׾�E�r���Z���Ů�)�f���XM����k��،�ײ$��^�5����,��������_:��eL��S[�*Y����>��m�K�yy�Ϋ'�����Pe�2�yV;�P�Y�;��lQ-^x5�������+�jx�]��N���R�:Y��(5Z�Y+u�V��A��hP.���JPuj��f;���G�Mc�R������SB����:�ʹ�UK\3 :��qɎ��][{���d	e�Z�(��_Bq�o��Ô�@c��>�����gg�َ; ��IC�Nh~4q�P�B~?]�.v-$�7�ʌMHңR�~�c� XT��ɶ靭�<|�=�\g�:D�� \�8M�ŵ. F�b����8O�^���[����Rl���&37N�_`�j����9��,�x~��P|n���о#Cԛ!c5�h��uȴ։��O�ܝ��Hq�]�iѭ��c\WnX�|:��`J��I9[	�"�>9��g��K7��9H�b��r0���o����5�ܰ21?��T��,�
U�r�ʲ�i��r���5U�5�z�т{��!���s��
�w�U'� �"R��o���:aS������Dʨ۸�A�i�>�Co���V�����1��<@g�=u�)n�-��E�̶���';�{�����Jg@�;���Sy�6t;Y��YSF��aM��]0�6bt�xa�p���A'ܔ��ү������zq,@}��~8�>��ǀ'#3��.`3"�o��bɓ�Ug���Uc�S���ֹ�`��ø�S�)�#�M����p�bo~Pv3F���8{��k�����ߩ����۠��Ҙ",G�Sq�B*��q�GU���v��;��t����#�˕%!g�⅖���ӉE�#����>x�LvcX�>���7�
D�6P(�p��wtX��Ό$�.#"�Q_Wq���d���A}�q�YTkcMQ�vg����"=�����NJ� d�,;��`ú��;?�o�'w���'mQ�c���_*ZC�+����B|W����tn9���b���:��Q*�]v�f��HS�F���k���F]%$y]�W�$ı���V�-��@������X�䨵<�|�Mh[��n��F�+q�B��h�}!�a@��!�^πm��:<��@����_C������t��z{�tX�Ϲ��bw���:� PW�{��*�Q�@L\i���1v*�rN