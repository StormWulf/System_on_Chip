XlxV64EB    40f8     dc0m$H1����4�DSAq̩����W4��$	��c>&���j݊���̪�u�6�}l&��t9$4�'0uf����`�&|k��^C�L�1pND�ɫ��X�d��n%[��	?b�I��>�(+�h$���4&>e5��6�:�I�]�
�� �o���z�1|W-s��^��(
]����������r� S�����	�.:v��b�Tu���e�^�=	�w�*��qQ�)��gN���5s�x��7g�>�/uG�$S��Êh��$�t@:QC�I�E5Ec�LۏQ�g�$�#��'_ݹ���a<.2�Ě�ʙE|d~:�t��\�6i�6�9�0��8��nx��f��ί^���}dA��1-�&=2�&x��.�D��g��$�4�T�#��đ��p�䵍\�A��Li�X�*D�u�ޥ=U�H���,�`�'�ħ��̘�С<�5���3�9	8�5*FsYr�|���H���2Q��"�%H��N��'q���OU.�!=�6`Ci2{��)%w�a쥵�s�[j����4ni�H ����=
���Q����!y�֩��C�q�{�P��DtJ�r->��֏�0t%��C{ ռ=h�(G�`��c��7�^.3˾�:�Fjh����~f���eH7(�/g6�u)
	(���N��jJs<��6�r��FJD�_�����7�K��g/�MlSP6nqb҆�,n�6w��QW�/`�\*�/H"�*�Q�T��� N�o!*�}z3A���w~(NH!���$ӟ]]����>"����������#�Yb=咻d�ӆ�VJ�ƨ�3SX��^.b.%�ͫY��߇K'ъ���	�z!ӥe�=� ���<����fm�>vNbG�W��'(s<6c�)iF{#�t���=������X�-Dt��*���Ul��z#�{ )�����z6U�@��>δ��< x\���0�Q8�p���gJ��#��'�����-���pp��w(#ez��iʪ j�6���y�d2n���>iA�g[�TY��✰)XL�s��"����	�H"�c��Lۙ(��*d��QL/-�g��j�3Y᪯�?t!�vu�D6?�є����`Y�Ģ��6\��M�v��������!M�c {Kq_?x����2<F%$�1(r�.�sK�(,E��_9��X�zIhH�w�snb�ν�y�5//�(�{(����\��&V���K�f���dU��4|o�&�]�a���^MN��A���ίf' SB?��9y�G�M�=���/���}t�ޕj�WP�=wn��s����F;��~@U�@�1�-m���C���������t��s#/S����A�x�]�`�s��Y�6ׂ~���(��0�E���
Pb��.��p#y9u�Ӽ(8���85υ��|p���Nw��En\veu��>�i�<��ƀkc���m�:����Ɯ<b�]B���l���5�$ {�h�pu� ��i�����)i4$�.nu���&b�5��`�{l똲6��P3�Xt�=��d��9�V�>��z<A�����us��M�L5������^����epq��x�)�sڸO	2����d<�o6kMytξ�j��� b�9���B̋H w�nv�en���0�ѵ���>�(q	ʋ���_��qYx'TA��q�ul7�eI��#6�H�,ջ�{��WϤF�s�)e��%~���P��~����)F-y�ǄDd�0�Z}�x��&�?�Q�Ծn �7Mت���E*�6=Dk���j.�A��,�G���I�PwM�n�8H�f�X�z��8����n(-�Z�DT`�q�m��c���CaZ�}������r1	�숟�BF�����P��M���5���&���tW�%e��	F�T�u�a;�9}B����tX���K�&���HA7[G��o�e�
k��˺��!�$y�:WL�iے��� [T���.H��D�w��^�}f�����lEN�m��i͞�n������w�I�Q�#�����	}�<w/�`�� �K�Ѷ�!��J*�r��z�n7!�r�����qE��MkT��Qm��ٴ�u9�$R�x��~�\�a�ON;P���_؃��j�^U(���~D6�=����BWXQ6xsΙxi�����Ԟs�i��NAw��{��PG�n,�{��aY��
���+������'����k�_���C���gd��+U��$Ÿ��mfȂ�v"�r�.Ȃ�&�w�?:mr��f������4�%l�]-n��^3S��{�?rWX����*���?)�.���&�Lf�k��Ú"��3����#�a�cȬTlm[�B0_�:'��A��������{�R�����Ҷ�L;R��}퍆F:<�>��3��r�:k[� ƠqW����`6`W��Ӕ�<���B���d�w@�zF����x��#�]d׹&i@���r.���e��.���ٓZ���(��P��#Y�~�����1�����x7:IR��PF��,B
�+�v^(����WNÕ��R��n�����j�"&B���z#m�ފ&�dF ˰��Gҙ/�$A�.U�i[�ݼ�;r�������m�E�`�)�OS��o�Ǥf�����=�v@�R',AA�#��Έ�gæK��+ȋ���.����h�{���4�RʗҴh��Kb��힑��p3uǉ��9�e>>��f�hL����eW��uVĥoW��������
��A ���Υ�FM��W���>onv�lπ�H����=Q-L� %8C'��<��;t6�ʀ{���z�P�r��������vdB,����t�X�*���%$�4���W�l��������k����2����},0̵��^c �q	�Z�ca cӧ��_��vw���t1���Opfe>��["�`��E�y\�q�#]<�O�������eADQ�̕���ϧ��H�SD�q'옼(���&�|�A���~���?�0F�3�ro� *��Cd��ANMEE�U6Ȥ\$��H'��"_��-~e0��x�������N�tB�:���˝h�++SK��=�)g9���<�as;���EJ�é�~	����X��i&��>Ǉ&�^�gY}��]ǰ��U������
_[)���Q����9�F>���˘&2��m�2a�=ǂ�m�}��$9#c��VM�e���$5rH.[U?b��ҡt�ĝ���̏ABN�1z�{!���X	�S肿�EP"�ixsl�DH$%ڰ	33�H~!�!��@�*�C<&؏��(+�`�4Ptk��ʛ������S�D��x�\l��$y�U�CU���l�2_W<;�WaX�/$:uv	����� ؎~�� ����G1��ʯ�s�)��*o����S��K#��i]eoC�󝺪��%���wPi�K�`_I7Q��=�uB��df��^S5@�HUw��ȱpq��L�í�()~Q�