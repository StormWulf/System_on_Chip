XlxV64EB    a70d    1bd0�5d����y��t�������߇47S>�nퟏ�� ��PDY�m����O9,_$��2�Ð˄0P,̇��P�ԔEb�{��q�84ɪ�?��Q���i*�#Đs(�V��`;Wz��@c[4\|4j���fA�`���q�k=~@FD���%@@���
-�Q�Q��&J�������oDk�]4v�uǗ�(vU'�qJV�N'�哠W8�J)�PN�7���+��/^�W�hTRE�4�Q�����$�>��8g��0�8���F�5h�rJ9֒-=� �S�����On�σ�3Oܺ��u�i?
G��M����vɯ��k�_( ��g��L+;t�m��|��_]0�Y�/̌���g������Ɖ�SFy�'����y�p��qU���'3�K�i����
o�����g���_�]�7��;�}?}�6��P��zi�15�v�uE���b[�B����?�o��ޭ�.N^�c������|C1,�ǶFS;�ok\��mz�8�.���ALb��@����
�S+�u����k���&7���7�b� P��t��'���S����S����1麖)�瞖WC�	
���w�t޿x(�>�P�1]���p|�}:'��cxL����@T��E���Q�X�ч�a)��=�څqV�>H�a�	�)R����g���J��i��q/�uDA~�{>xa4��m.�GQ?�EEp[J�/�-�7#Ӌ�tИ�=�&���+E�x��G�s@[��pji��Kk�k ;[>��=�G��QN���w�{�`_��1�P�{�([SO��1ǎ#p������\���8��E��H��:>Zk%>�`E������Y�k�9��אT���Xߤ���f�}�qŰ��AxW�c�J$��h��-{r��i�mws:������P�B���p=X�>=�8��IR$���y9��2䌂%!3��D�et�/��Ұ|q�ع���ʠtgj.J[x>�H���dR�O����Jj�-:f�+-�}u� �"�WC���qG��R�������f��� pmؗ>�����$����>U�L4�Ȅc���}q^���Li��L�}��bhb@U��I)��4`p�b�8b� ��&�͏Hh�H{01=|����4���*�_���HL�/?1��lE�� ��p=~*gX���VL��[�`��o�I�����7R��Ѯ����ut=PlӒ�Έ����\� &�i�*��2V�;`2���`���S�d�!���z'�?���qT��n��c��m�D�FzQB�r�,i�e�
�����2��+�s<��b����Uѩ��ʪ��/z�X��ς���PL������>DV+�a�ْ�WxZ�*=X�0m��(/O#�y����U�u��	1�f��<�,�����{��5S����s�� q��l�,�x[���!����K��{�E����5I�y��-�L���3F��w�	a�9$�}�ف8%�4�3uC���5�p�pzi�p��N)��fYs�#�C�%��pjOP�oK�Ï$��H���$lۂ&����O|��B%~2/zp�����h�{6N�>���(����k��9S)!��tm��X��.`	���h�8��.!o ���8|
jXgt�N��������øg�ch9~�Mz���M��$��H��߹����0�#�sG�䕣�KR��0H-��[�V7$m���BD�d6){R�G��=�6'	�#�"LL�6��8��ػ��k ���: �<o��!�s� ��0v6�l���%�3���@/�H:,�n��a8vSA�����іS�T`��u�徒��j��/�B��(�晔��h��� �K}�n�{��2��D
~Z	)0�x=-W
�o+�@��o��ŉ�'qAl'���4���K��R��1G��b����W�er"މ�Y�� zͧ�iz�*����Y?ӻEg��$-��,�(���t!v% }���	b�1�!���#��J<¹"�>3�hW��;!g��2�>��3�	(#��s�j뚜��kle�-f��	���R�i)T��b]��(n�8���6��!�t��Rd�����oN������J�&�����Qm�Lsh'ϲ�3�a�#��r<5�'d ���AaoHC(ۗ8�F��T��J�V��ܷ�$�����A�0j[�I:�{�M����w�t���F�D��g&y�_zoKL� �,_�R�	��DI��B��'�����BR�U'�&��Q�D�	�+�V�^�[yx���V�R �:����	hHY�hh'qb���_�{ܿ��oW�U^�׎���*���H_)_��ղΘ���&}��b��a���V	�	6��"H��:�yܒ�w�RQ:�x#���)ʪA��@Y��F��b�4����kdSPO~�[�u�J
-*�G3�(X�Hn���(�6�b��j�MV�7��|4D矈�oU7��0�<ӘiD�m6�S0XT�K:J*�f�с�����d���Rn$�:��8�M'*���B��]�%�&n�Zg�V�P_��h�n���c(`8�V��r�����n9Ti���B�lyH,�!gJP�K	C�|���&��Ѩg�b�|����o���$�7��B��]�)dՂd�d��-ҙz9WK:�=�QT����߷��ENt��x4�=r�m(��'�o14��\ȾU��EJ{�
����[��$���;��<?&�.��e��ϥ�6v����� AX$	
��AM��pú3-Mqu����#~�r��v��EE���>=��=�h���ǿ0r��&eC�0��?��`�R��9�TVp �j�3�*�8�9��`@��'9����� 0I���$�L��pD��"�r*��!��ʴ%Ýč@k#:����r���FC� �z�9�]�Qi��1S�_q\V�]gX+h�L�u!�/�h:�|(�
ݠ%4��!�]��zw�*jIJ��D^�gi�_���(3�[�]��`�w�P�m1.i11������b�ђz#jn3���Ȍ�m\ �b��W��>�N���z=RŚv�=��WU�����HL�VNz��_HfL{�w��|hv�ޝ���ձ�%�p���$@��gi`�0Q�s}����d@y��0o|hn�"�-<|��c�Ah���%\��&kB)�m��S�C=n/*��6y���TH^�ve����E��n�̩��[�aw�W��%~~ՃN���.�P�y�D�^�m 1�E���y�A5!}8�9��U���3�3�#�^��(��3�ȋ�䣰?�B
f���j������K2`��!��'fŏ���s@Nm3>ڃ=��3�G��$�8��>��[EK�9\f:$��|3���ߥʆԝ}1�j��
�����L��e���\7��sX��{�oፋ���m�U�8f|��Xg��S`����"��a�$��k2�,��=�  �b��� �b_�%8�D��mf�l$��-o7��o��Q��h�?����ٵ0��\rj�����v��0��L�л�܊#v�]��l졚��,0^�+�b3й��M��=d
�2~�����/tk�{S2Y�VJ{Lcu����(�B�W�Ħՠܿr��x)���q �g~�T��3���¨������#P�d����=x\�S�j������A!�+0�OK�����Ȕ޽�͸�J��?0��P�V^��S}]�p�B/��(C�W⹡�v�!���1���K��mNN�AK�UN�ks��HӼ>ki�Ytڼ��§Q��4�3���b��[T.�݅#��.�F/�sǋ
Va��!l�L/����s�zq��M�ᵀ-�B������/�i�9�N(Ì %��W=�2���G%�<��/�ǷA��!-ڈ˒��/��/%_P;2��F�*+
�l�6Y>�	�J��D�e�8��#�B�qNp�4N:l�+��l�{7����>�
U�}e�mp�}}�Z���sz�n��	�σ,܋�R��X=�"�&Dg	8�\��vM|/M��d��տkCy����Qp#,�[<d��4��~�c�?꼢]�
���4���VDL�-��
����0�B���f�;��N<�n�����!�q;땟�&3.�1[9�_�}&���p\����a^���N�r ����b�Kn(��`(�E ��� �v�i9�����媩˱
��$iT�c�o���I�u���Ck$���N{�$zq���QL��Z}���mt��f�C�H��ۖ��]���:$�m�]�K���ȃ�~�TxWDv+�J�S]j+<�]A���@���rP���?^�ގ���K{��1#x%��lX'���.P����Ʀ��uaS���3��U��O�K	<O�_��P��Hlo�k�q�ԩq��i�z�m"�M�ܖkw�w�|7���\u�q~w�֒CC��E4��>[8`�o-�n|��Лe^�+PN��ξlo+�C�����\[�i����{H��+D,"����EF���P�5/�$n��4�XX��&
������vc{�'���z���,��5��1r,)I�^i�ǎ	��6x����-�F�RJ���h'e�^P��
��0�.G�����-\@�d�4���i���&U;w�vls��*ds������RT�Ih,����X|�[�ο
J8��*w�5�c)I@/�FV47ĉ��lwu�rʍD(�k!L^�k��|=�o�Xv�cb�z��E(.+XRN����:�{2=g'2�ϊɗ�ŷ2�����
��r�����V�
f�R�xT�U���Ӗ��KTܨe��K^(���V�=}�t��i���$���#��d!�\_}�\Sb5��?]^݅aH�k8;-���
Noor�^��:2L��T���9���:^ �@3\^^ĝ�A��jK��	ۋ���b��ң�x��W�Y^�����t��$o�������!N�|�M��x����ҡ]&����q�K�@D@mַ��y6x�
x%�� ���@�N\Pr"w�h��	"z{�ȟ1����� �R����˪�B�G�Ph��<7�ސ�ʔ{�|��"���n�����5��O�$=RY���K=����x��+�����IɆVdˁʨ��Z������H�/E��!�E.��I[��{�p���[cç�d�n��fZr�
�VBJ��?�uһ�t��e^�~�r_�t�� ���ڛ�٫����������%�) � lo�����C��w7'��b"�c�23�0la���.P03*b?�Wm8"��d�Ml,nk�@��8(8&O��7vȈ{�Pv�TT ���&�rtN�-SZk��*���(Q~۱,HͿd�ߠ���F�Fx�r��C���y��#%5�m*(��x�t����(`'4e�`N9�͉�m��a�}��D���E��Q-��d���ڭ�:Ȁ�7D~��`�j����h���]װT��n2�(���d�v�E��Qx�L;"B����\���4Ԙ�$�h놩τ��Yt@ӷUF���Uu�{�.P��?N�b�Y�W��&Ju��veg�b߹��C����A�q��ܪ���z/�:�b��#9h�*�~o��'���K<Āb�#�Z�����PnZS1���ft��ȶ8�m*Y�<��ƍ�:Tp��">a�F\e,�~�t���(	��fxi��f�qh�	{�Z֚�Q�agו�n9|C�߲��!@�JHa�����VWT\�`����=�n.�*!2+�(�� �<TԦ�1Ey�#�U~��(K�xa�yR�8
�WI[���WZ��t��Z�YS�񨐒�W?O[-O�v@����C�*8�3-���QY��XgN��LiS4Ҵ��ٍL�b�nc�;c2��@)������L�AP@��<_
��oRw\.�=�%�&��S��[��Y��(���D�w�A��h����R��D���9X���ĢD�Qv	��X^*	bz�Q/�F��
X[hT�J�b@5���!�,�f�0_�`��r���U�娦�S#���} �f�/DX�(/����`�#T�p� +����$hQ<i���B~Z/UU�Ry��-��2u��$�@��f�58T76ft����/�]+#��HB�o)����xG������#F�1=�f�����Xv����8d������R��0U1x���BQx'��=VD�	:H��@݅n�i�}�#���_��v����Z��D�<�_�=��B�1��8,y��&
6�5@�Tvy�\�������M��'c#�O mn'w2Rh�A�)I�<���.���[$�e��k�Ӹ�Y�&3�@=:?DGﺢII�؅��p�Y��9�'7牽z@ޤ�@y���k��ה��m;����u�I��H��=N��u������ݷ5*u�'���o��i9J0b2+(�J���)�ff�O*UL��ۆ���-���"��hiBUfeTa�,W��aټư�B�ߣ�iv���������(.�-r�U݇*�gfJA��x��/剖��ڪ�H>c���]��3�bg�����Y����Ѓ9`���ϲh��E"�`�����X0R��4�!���=v/��0+�@'k�?������7"�.�I���ǆ�Q3�`����ns-�˺�CQ�5��Rm��յ�=`���"-�h������fb���e{�z��a�\�t�c�ߣپ���>QGO�#q��N�W�S^�{�2r�e� �̃ѐ�E,.��������������\���Ł(����i��p��.�#K�3,���D�9/8���� ����i6�2��aS��>)?�m�U3����h+��c�����L����`��d���"]I�T��A�8:��W�����K�f��M3�i8r�VԂ\�F~,E���cq
t�Gw3	K=7)wK7���ڮpΞ�ű�/i���Cv|�����hɅ�;���O$<�N�����~X�(D7��x�3�� ����6���ԟ��