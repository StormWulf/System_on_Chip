XlxV64EB    3a22     ff0����XA��_�v<r����jg� �q�1)�>�YN��x� +.'m0��{$֦A������#��P�o������tF�]}����x�T������������y���S��.VT !�a�&7�����[����u���H8�_&D;�ņ��Ť�fO
��D Ԉǽ���N}ʫM2��C=�:�x���T$��mM�T}$*��r4Uy[��˛n�\n�`)π����ōIp�î��@fg3���1�CF�p����G.�22�ͮ��M��+��x}���\���B�m1PS9�9>{�)#���χe��m{��3XJ�EdZ�O�	��7��~��d�5k0-k҃F����O#v��4��&;#��zo(�����@u@8�<`eT/���Eƾ/�d0�����"���mS�B�W�s�o���TbRp��;��4�?2F�7a�58C`�	��{ş��73��S�{0�6��w}��,]-�n��Gΐ;���x�R�!�\�uǗb��_:Hl�o�Ķ���}�W����}�s|#D�����"\4D�.M��FV��[�6W$.�Nt�r8��I2����0���S���|��Z�)�I��C�G�)~yl/��Ay��W�G��J��U7�����n܆��~�{%C ,��A$0��,���I�M���i�H嫷Y�/,*G�Ñ#��/����@0,'�3�1���Ui� [�D�o�s��`+1�l��XE ���}�8�{��c��)6�)��"�[w�~u���T�k�� ��'nb����y���!!�"�r^�9�Z׉�{�J�xm_�I��*�ju�����m&�D�<�@m���_YZ��xpZ������4NÕot2֕�qZ󜤑�c���;�3<}��
<Fm�
$Õ�8w8!|���	A`2^��)F�<,���n��u��$��Ӽ=yW����MPj
k�D��-��姨D�A�� r��Md����c���b9�Fl���M�G{�Hީ+4�k���D�3�p�:��)½��qր�7��Q��4g�6���Cw��:�K��Uh�������}���@#�֨��@|Y�L����F~�������*�ɫg�n
5�}�X迵Fo��j��&�����9����}@��h+S3�~��؁��)^�{4|�t;�>.A
(߅����RЛ���{�)�˺�ʉ`ks$��O�Q)w��Y��οQ!��)-K�	6��ǿ�\���S9��I���5�S���	�b�a1�7�$�.) hC�W�"QrN6d�r��j��	%�y��G�X�]"o"r�Ӕ��=+c%�K��}�?#`ҷ���v�k^�-u����m�['��/�׬��M�e2.9)]{Xш�'Z�|��g�<-'���Y~ofO���pT�F!:�]{�Z�w�����{R1�\�u�A򩂆8:�ÑT�!L�=���+y�qm;�CF8Wضē�_�TB�<uΈ ��E�� ��!FtH��� g彆2yې<�z
F���s�#���K��?��F�M����cm�1���~����p���W�&�\o�ǘf���h'UȰ�R+0Qxf�U��t�HxA��
;\aj�j+�f>?$�p�]N�_f����igz<_�h�}�I�����^���m�T�@�ʅ BO#��:�נ@oU5��#N�@�	5\�����^A%X��%�M5l"v�/��ۦ��TO��]f��\¦�oQ#�#���}��tr���^M1�C���&'+��u�bO�J����H���# �x�(B��D!jCx�b1��u���s</��`@i䌰��S-���T&��PT㦹s�q�e�ɰ��Ò�;ؿ<�]���8vBK��e'�O����� @ѺzoF �n̜�ύ������z��s��\���3�� >?u�p�:�`9f���^|떭�ޙ2��������Cd˚ugvA��?w�;;̍�m}��_�!�9�h�o7��h:��8p��+��`ł��� ��I+[[�f�m)��n�������U������`G��V�LuE{��D�m�7��{͓HY��w��F�q.���ߘ#̩`�6MÊ����]�F�i��ؓpSC��-Hdv�l�������Ʉ��a��������b�E=2����m2ʼ�.����7�,V&+���8�y��+�NTy�{$c��i��@�6�/�(Y�ע�yہQ@�D �@uy����Y8��D�u9]P�t����! ,���Ge*����	׉H� *iQ��U0ؚc�A�p$�΃8~��Atp���赓?3��@�[R�j�)�\]̝\����c�v��ʹ�~��?���P�r;��ew"��g�c����w���܃���W�4@���g�`��/��:�������m��hS�1i.v���w�~R`z���5����n�'���1:��N����T�ZĬm}����`Qo�67I�m�Ϯ�OI��I���q\�t_�;nƑ����}�%ʱ�כW����3�fU_������=Kb?2}�B+3x0G˫���[hV�R��0�҃�������7���P���1��N��NY�v!�V�����ׅ��!�P0���;�_ܣ����j��ۤG���6���B"��u�x�Ʈ��y�"{#э>��?���,]ϬR��%��@��%����-)���],��\j.�~$�B��\=��!r�Sc�+8�H�R��V=�d:\d���++��K�V��CŽZG��M���j^�FM��10���j�ʶ��,�S��x�zemE1:��sL4񁺛yR�,$h�^<����?@�%�̷�)�lES�+ń-6���U�|k�����,��k5X�@���y���|p�pB�H]3�H�]�~��Y.�{ͯ��:a{��g5񳔸�z���pY��q��`<�=����ఖO��/����?����8�<��~� <c��p�JYwJ�X�"�X��Ġ�ն�y�Pʐ�L�A��|.ȹI�Ak�k����U�G��{��3�e��M��� ���� ��׫(�U�������5Q��֦P��qF��R����]}KV�6���"gb����{���n:�e���2FS���hhc8���;(�լn��k�+��m�ϧ,�(Y��6?z�NQ�g~9���a����0��CO6y�o��w�-<����0P��8�| ���@�YG ��N��M�P��1�x1�
��8�tڧ��w&@8��N3�˂����Do�%�sc7����%���G*�]�NVh]+�DU�!OY�:=����AqF�1F��%劇^.Γ=�~+ %��Rk��R2׫0��^$0[�4����N:9��:���:D�����8�D}b����k��f�3
�K�$���j�4�Q�����!߹�������Φ�@gNJ'e�E$�m���He�)l���>͎<>+��h�~�""�@2��Z��KFΓ��uZ1�L�]џ�7�:��Qwc�썌F���h�jzx���Q�O	��5�����8�l�$P�i{n��5�@�)p��0�߳zV+�(���� ���	���..	�A��hG� N^��R������蛀��;��5Weod3��z:�$�����D  ����c�gG���sn�=n�8��Z��.�Bn>$��]b����b�T�y�D�:�`q���A�}�:�+�����/>����ʭǎ���}�V\C��l�Z�������Z;H���wX�m��ʓ H���LԷ�A)xb;��N�@�gA%g���7Zl'z�Ѹ�Լ����8�T!�=ϽHy�:�Z{���?���v��I���0��s!��9(�Kaf��h���
֖J�E;7�0��t�v,8U&�fʇ!��/+�Ȅ,�'L�8�2�W�䰒W?�Òci@dt��mbX�3�=�!2�$Oٳ�3�W��W4�ihZ��ٔ�)�|	�� mעT��� ^Y�lD��mq�_,m�On�	��=	��_ۧ�˿�)"�9