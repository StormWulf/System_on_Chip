XlxV64EB    1945     9b0�F;�\""K������ɎL�n~�z�Z�B!�ͫe]�h�s��_%0=�ߔ	~��'Ѿ��sMf��d���jG��Ӵ�mD��Kk
0Ц@��
���}?���TU�4��%���Ws���(��D��;� ���ةYpK�0���u<!{1LA��d|} �M�%�W��r�L�l�p��|���u3TG��* v���L��e�� ��L@a���A����e��o�����+q����6��h�;��2um����*�a�K�����}�%��d����ώ�]
y%#O'-5P�q�h'�(��z�k�8�5� �;z�;^��_��l���81;o,�\c�ԅ�X!����D脋��R�U�2������G�fs���Ҕ�<1[�8�k��TҰ�S�Y���9T��3@"*>Ϭ��"F�6�D3v^_w�yU��d8�&���|b�0�_�.:le�X������t���~�ֵ�֥���S����7��k��NZ�"b՗��"�z3vE<bk�?�����_!%���K$���1W�n+��}��p'9������/�U���s����Ƭ~Y�㥡�h���cZ���K�L��s8{P�$O��p�t�1�3�<)�T9{�T"z
���?�v`fFL�f�z�;-L��s�{A.z���O��
n�(dA'��fo��ǚF�N��J�M
j�ֲ%�^�c�:�	��U���;��nq�h��0��-&���,�<2�p�#m	u�m]	�2������39M�� `���-V���v.���ϛ=�{~�'>���Q�?�dg������3w�&��u2$��˱}�D&�me�ʌi��#���?>�'���G3����Tb����O���ѵCQ	I#�>�|������J����,�>�yؘ����"�m�'�� � U�}��Z��&�&f:���q���uw}S��V�%g����,��)J�j�^
n[<5��M�ߠ׶��tKvY㿷D_q��*�0:B(�Ȣ�20RZsW�������b����R%�i����d�w��K_d��~�]��p2�Т��9�`ҙ��P1h��?��J���;��7\�X�����CZy��ꩂ↤`�<GEP�\�N��%d��M����N�ޫ�O ���Wn3���nm�[$tb�+2�˫���<�x��O�Tus'4%�����kh�I&5������
�g	�2�^z`!�;n��F�	�1�|/ծջ���.��P4��M9��w$>����	z�[I����^�E`W^�oR�^�l�W��zm�1�}�1Ґ��������|�c&�V�k4��.<��Ȋ_�i���6�̩�aͤ
�$��,ŷ��Vv��� �8E�/Ɇ�a�Ek!���6g��~m8�6����nS~�'Є)>�'[�d�(���fa[
���\A��j4�?M۵�f�Q!M��E�em�u���-���?�r�`�:f����գB�M��j���;���aJo��[$��w�<.��7>!"u�;a��M�FK0K��^�|`
�W;ƾ������pl�����D�Z�&��
zmD�:��߹���I���O�2yے�;�ӎ*ZE��r�>����#�t��WwQ#���QM�y�2~I{ՄJ*I�f�\Ap�i耥���%�w⍄���g�E%w9c��,zA��9�@��Z'vyZ�ҎY=��L�;-1�,��z�	�����9�_{ս�J��p���|�-�B����W}9�/�-�I��gЭ�������0��U��̅�fq�5��[3�8c�6��xp1��I��mӝ}Hd�ژ{���j}S�)���Ԗ[���h���� 5DOl��J/�3�ϥ#Դ����]$��w�c��H��3ΐp�*3�|U2�������_�Ŕ�hk� ?�Ϡ1��d9�1�Ɛ86��i
�S�,���S%?NZ5Ԓ�i�<�t���B��� 3� �|�1��qX�͘c���7=��k�Q��e\����%�������/MV|�%X���8xZX�|�ts�|�1Y���K�( �@�j�Y�B67�f�W&J*q�W_޼��_8�1|<r�m��@��ď��
q�(kU>�����
�u{��Q┍���,���u㷅��5�����P���.,���0����dV$ʇ�1�T���Ç>Zi�B󨽯�o�5i���X����.b�0�	p�T��6�|���T���p�t�6�!dL5ƴ�j�a��>�-X����c��N��?��I��t�Dv�|>�^�S�I@r��n���p\b�0��*�ګ��w�OWc|J
m���f�-���fh���,@�tT�!*���6�m��� ۑlZ/<@ }7I�w��s?�4E��� ngz���z��Ft�B���]���cYu��
�@A%�p����ub���k�ˬ0q����' ��_�-j�&3