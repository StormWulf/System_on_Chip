XlxV64EB    163e     870�����:L���Ν�b�W�'��K�< �`V��b�C�h�8�}ky#�Ԥq��G���ߟe#l���M�Up�����6%\;�I�dff L#^\���fm]E�7W*{a{AV\�a���jFvι���D�0 �ܖ���-/���N,ę�R�QUi��L��}�Ĭb@��ɚ@����>��SBY"r����S@iQ�����7`3�7n���p��|д;I;A^HvP3�n<$	��ݾ={v���4T���s�䵼�4޹��G�p!Z��4�Y3��!8�M:�9��4>�	��DZ�x�.���D��{���iu�s2�21ǎԪ�7%�9�"�n��ic`�%�B1]�{
��;թK�mY�(f� B��/��s}�0����pSt/:R߹:��� !ad��m����(M쐵f`���7���+�S kY^	�A��B��z6��p��īЄ�^k��y����4zʒ������B�=�F��fK��Ŷ�ݻ���+&���Lo�R�`f����>ܮ܉`���{�aAha�(���|�!I�h�`�@�y�?�|���L�ʆI3�3�����(������K�h,��Y���3�tJ��8~����H�����ݔ)����k��n��59g�\Y�bm~
	��J&���#0���.6-F�A����	ؘA�H	���Y2���� ��Q|ȷ®���?��zb.����H|�@�t������Y���2̨)�����]GC�%��5NA"���N}����d����)���͎���'�.���v�Q��I��,�}g"�h}�c������|�L����M��2��#�7# B��r�)l>K���ڄ �j��LQ�.|�� ���������R�p.��MA��b���M���5�9���g粇U?������2�_�_pz<��Zuڪt����%��1.�*5���g��1��h��=ŏ�widV���0���Ҡ��N��T,^��7���}�����D��{���0Q�tx��г��p�������
��!��]�ㅶ;�ffB�[���IjqU9'� 
6@ؑ\p�kzmۓ��T���y*ˢ�D�]�.7��O����e���O���Y�۲,׌}�I�=��/]�Z=���;����6���yn��6K]͇��AJ�ξ�����#>3cb��PT_��dak��:��|���YKz]��t��zH�|�K��y��I�Ѣlц|i��IfgW��s��U�9��Ȓ�e̱���i�{g�(�X����i�j�Z.���NK��6�R�ۈ��W�~Y`������\H/	�R��<����m@|�ɍS���C@2�]�}"�-���w3��on)��ߢk��٧��7ФDɞ��f_7��I���m����:yRI��ZVؐ^���r�d��� �W�G��F�����?�OwV��u������S7������(�1ޙ>�/i6&N�$�����7���C�[�S-")��#c�Ļu�t���RP�������L?�wqy`��J>\�[�P�S03f��0������PE�[8��)�E���D滙�������*%����n�Sg&����[��I��p�*
�/=pM��tJ�?�����k�>F/dabgx83�e2.q��`�Nƫ�^�"��+*10��B��ŽGe�*n��a�ro�?K��U��Ƚ�~��~�jN($����Y�6�5���T�0��\h�3���]S�t�`�#k��陂.��\e�=�S�B�6�hu\ҟ>r�HQ��qˉ�ON�yS���@�������>�, -�um��)�[��r�U
��)1�D��ڢ?x&�ƙ�&�Z�	��������/,�!يȋ��o*g̽��>����U*Ɗ>�J����M�ufd7�������BRҨ���$�Q� �����V��*�7�����Y�|��aBy��_��\��="�:q�` Nk�߻i��v�ߊA��ve��~�����o M�� �]��^(�K�n�p�!�O��i_��za�R[V��L v�ʁB��҂����D�����������4���8�K��\���Җi�&n�]W�����rF��W���V�V6��[