XlxV64EB    fa00    2b20?0��DR9eB(j�-��������/�R�N]�_D��j"tgJ��2����cʴ��Nn.ɣH��� �Ē��o��E�u=~b/^���!'|�6�>�x�ԧzg�5��o�F��I�S��3�3/�7<���b�}Nx��>Go��{����,\�����6qa�2>~Qך����vD��_��3�{�}.k.�_$�=ǈ��|}ûc��(W�u�&�.uS�V5�]���(}qz��s>3+�R�Y�@�\/�%�_>Qfh�5��F��6�����Z"0[s����K�2#����kƎ�p���0C܁���j��Q�������L$D7y����Y�cN-�Hn�ۜ�b�k_�z�.Ϫ���a����>#"W�$��L3H��f�F����3)�]��X��S ���Nj̭�x�)g�(���{B鸐��[xk=�x�'��v�7shː}]����v� �,Z��
� e�mp+�
�S �:��\�N�&`^x���b]Z�o�d����kP�^����n���(�-�����?�.#�˧�E���Ձw���8$4S`N`g�&a}�;��Q/��P%����xD�d��`��I*�	�?�s"_�����B�������‸���y�������?�� ��{?�*�CƤ�f@C�ưɊ�m�2��˫M��A��tg��!����J}�w���=g�U�E�2�cX.T���P�����]�Lw�O���v�`����t=���@��^��% �����Rlk׏��V�rlP���g���.�5�x&��̋�H X��黡l�X�@m�Vp����#'*��Jfٲ��UW8�
��3fH�<���K��\2������2��TKk3���w�h;{��>��I̢�+':�7����xK��
G7��{�`�3���m��I��$�c�	������-�Z�AP�%����ԓsH�+�J���7[��ʦ*��T
r <��5��������M�'L��*�J���>�����Q簾v�s;cGR$�����D���i��,����B�Qm��a�8T�15Ag$�5{_ ]�w.-���	�xJZ�����)4�����*�G5��W;T�th8�KLG=l�U�+��"p���c�,�k��"n��tT�=tܯ��7*��Y�R��m�C��� xƕ-���ρ=4��λ2(�����VA�u�e�^+��R�g����Q:� �O28a�sEEԴ���t3�۔�Qĺ��Բ,4=w%8�Nqs�)JDiR�8t�-�N	{8.��|$�M�4���+�f���2�_q�����_����9���Wf�gr;��3Ӡ���.q�]Je� (��Q�>2m"J�&��i�
W�߇T0w�ի(��~����Qp@0�G�D��V����5ޠ��*��59��%߾A�Dh���)�K#_	J��5G�3���X�,�v��h�ı���;7w���R�8�
5Mź-��3Gr�|��4��_\�H�.��{V�[�=�:EW��Ӽ��P��¡>b�"�>����U�K?���c���Mv�$���#SY���h��5�9P�%�ۍ���
Jj"6�	�za�8�If���]O��4N+oے��F}8�)#֯�n�)�n�;;A\"�O�:�o���W�n�N�
���'��Z�nL�#�rN���`�Eq�*1G��U�AL@�W�:����5�n�����~��`���K�B��= [r����QF&�D9[���/�ΘZ��\��L7� �Y$h�=�-���yCު&&X���ΣY/ޜ4�p�������MfI��2���������d~�Ԣq�PĿ�L��+��
=����_jq���1���UFR��8;����F��͎��f��g{�w}rH�Z��J�\wbL~¿�*@i�[t�*+�3���?h���|   >�hbp(��1�m*���B��`v����~�si�	�����]e·2�,�����<��ԘO��WV�.R#>�_�۰hL-�4�Jg�͛���b�1� �O<08�M� ^�A�l��q�{���g��6�!S����h ��S�&��tmu���Y��M�}j%2�`N�K�@_�v�b@Ri�I��̟B� ��	?��J=���Ɓ��-�RsV�g�QS��.�B/�R�y7+�Xpj-<>�\�tD��(v�Ǡ���ܠw��n�W�z�x$$N��"t����tZ��L����ǁ�anᦇ�|�_�	�,8'����Zi�����$\V���z��B+a�E��!v+m�5$	k_���cuG֗��Y��ٶ���Ǡ���ןML��s�T36D�������Vx� ޽���@֮X[Z��^�|_f�����4�w����;�i�vh)/�G1���]�Ҋ5�r4�a< �
@[�j��;A�����G�i��9��V-֠w���l1�]kAm��Td3�h'R�ͬ*"����ۗ������6�@���(�������M&�fTD����ɜoF��2�y�;�4ͨs�v��u�"�S�Ｊ�{-)�y�K�&QR��5�#�a܅��3 ښ��A�Ƣ�)�E�fV-��b�ꊣB��]x �+6=�������<�����mz� �p�0�dS�F=0k[����5r���v������mCv�ʎ�NN:-�<$�-xxT�Y	jh����x���,�Ҧb��X�oxz8�2烉�:A���ͅCk�-�^�$a�;��v%o�цߞN9`���3�рs`T� �X����xFk���4�X���D��k�ӽ`dį@#���*������w���T+T�!�6pU�v���^�������?��F)w��.J>��-)�E݈��iˌd�2�d5;�p���4�Y�
��^�t%���<�ȇ����l]RQo�V.嗴�GVB-
��8L��e�iԍ]�����jo��ۮ�6�h�x}�:�t;�7�����S�S�������_�k]>�x�AK'KY9W&���"X�9����|�\����R�<���k�hjl9�"�_�:m>Pŭ�v�jG�i���Τ��/��h���o{�+\��/��S��Yj8��f`�8|�,)�[D�6R��Ya��Hy������7�{�t]Z�^38X7�	�����1L+T[@��r���EQ��}��w �҇[}�^�$ͮ���ʥ��s�_�-kf
F�Bg-յy��j�7
J!�!��-�)	iڟ�VXJW��\}Ȯ����#2Z�J͈�o,f7l��.+>>�BݐL5Z�kw
-��g�c Ԫ �h�;��)�%�x���b*�u9�x��Yʈ&��l����s�D�Q["f����>Ez2u�}Zd��{b�"�ìn䞲��t2W�����A7�������9摴�"OJ�OJ$<bA�SY,ލ����v���)+~{���d�}(U�Ņ���7^�v�|�7E�qϯ���H���
�xc �MmB%w�Ĥ���'�����_Yeq����o$���������x���5�xYQLA ��G$�0~_�p��s��Q����-xl'NBnU�zb�	3e����F��1~ए�C��y@�)O�cr8���y��E�i#S"ȴ,Hu-ޢ�� �%��Q��6��aG"j+�[n��]~��h�"֝赑����%)t��h����I��I�t�$������6<�8d�iO���X��i������\:�fՔE����j�D廉e�GRP�VjPn���>?Qb �0`�!%�6��l��#�?&}+�q�Z��S�#����7�c�;V{�E�m����&?�G��  q=�
W9��/����H|�NB���	�R�]�qU�%;G	�d�F���,u{TU����Y��tu��l�>�@,��CXM�2֗�G�퉱z�
���f�y����8y�I����q������g�M:
"ԙ��7���#^���� ��)u�85��l`�
�B�;m/� X�h�I%���=�rGW<���aF��/]�D�{x�|(^p%�̝d9qBc���
)�j��\r۩��awQ�q���V���̼���LJ���v����S�%ǦS2s"�Qux��FM�m$�{��ݖ�5V����O'%�"/�� �r�I���hJtl��8����M]I1�F揽I����8��`��ڥ��p����,$+\9�z�L	�uK��
��n.�U"�X82@��!;��P���nl����)���̵*r�����y�T��WG�8k�g��ʣ�R�*�4�)W�}PMf]� [33w���X	Δы)�W�Q>�zx���g7*��\�O%� i�푎�d��h&"ӷ^{�H6R�9��jN� �d�W��A������zm���/���xى���W���jRt �FؿM���z��������t�������p��vb(bq������x���=k����iK�3VxR�7ۄ�dosH^U�*�)}<̘���r�{���1qvc���� �^��5�{�x{�7�0�%qS�!��x�D=��IG�ғn=nB��4��bis�
��`R7\�s���?�BR{&T%5`������:Hn=ɤ�6l ((��ΪC�Ӵ_�<\�����
g��b��r2At�?;�L!��M0G���>��o���@G�b"������m��«H�����tUUJ |J�Ђ���;�!��"��X�Tnֲ��w�Е�(�℥eE�E�E�m&�L+s~kD�9��&���/��_m�1t��a����M��@Tf`W\�-��.���b  eyU#�}�Gp��ox*�j:��!�sOsd�]��[����G�!�ywU�^���|wxQ�H
b���ϦR ��9I J����΃ԇ
�|m�4��cH�8�֗��V̼���-��/�/��AOv�n�h�:*�������FS/'������{c�����F��T��K�_N��L:��x	��9�5�aqL�]9wbc/W_��_kA�*����*Jo/����y�ae!Kp�ݙ����� �}X�^�$7k~ɘ�{��i���Y��N1^&Ӛ�O�&�V_����ژ_t��d4��[_J�I*�W使V��w�u��d��oۑ��E�EG�Oq$�F`[�
��NȚhxl���(�k[T�\]�W�9Q`�S��:\wa�Z�R`ظ�[1�7r��Ho9C�ݫK�+����=�1;efv@�r���yf����c�Ib���S��B�4����� ������8̞�q���Qڦ2�Z�3�`,�=n�?���7���/�#�˅󆏮R������*��ѲY��n�!�y���=p���Rmŵ�+i��V|�ɕ�]EN���pqc㨖~bt����Y���"&�O _��[y����w���D�|�H�S���
?�������^������4��V�֠;�s(�Ӥ�9���Zٙbq�}�%�%ZG�k��x����=�Tuӊ!g��h��=�lre�؍k$���<}"�Yԅ�qŦ�݅iΞ]GH~ �=˥��z2&n�4���g��@N T��ƹ0/"L�6���i��P=Ӛ�ss��HT�B��P8]:�[�I��a�I��
��1��c:Fgf�v篤tҔ����ϭ8��|��5n�f��D��_���?���l�kl��.	��(Z���j�~���ASH���wSW��"w^_�e�T57?3�"��Z1_���)�b��9�f�t�!�~+ǖV%/EV�8Ӷ����2(e���A���hU�Y>��9P�	2��6�����Wj��Z��ꚻTD0��bO��}��h���4�<v�>��Q�Q�  �K�#629e)N���O���3�<15I����^�k����S�(�u���A%V��2<�L�fIhq�����9����V+I�	(�w�eN@p��j߱�n���3+�����&��/�+�3�uE��HO]��I�K/Ͱu�1����I�
Vj�a-5�D@��t>�[mc_��tP�w(�c9q��.`\�+��Hu����?t<�鍎���5��:����i��^�+��Ê���Ϩ%9�h�E���Ƹ��EQ�,{�+�������e1�'Pn��ˎFm4�@��~7J��"�F�13�f��B;.5�&I�_����a�Xޭ U�� �[�R�tE���j�q��qگ. �g>5K�ί��.'F��Ab����L�z����v�G錿��e#w1��N'O,[7C�z�	�;��d�`�u�2����L?�(��ӑ�i_L���h�G���(`lx�s�?��7�y�_j�fͳ���W�V"6v�\#����fΘ��"��h[�~*����{|:7��22�V�da�Gm�%�?ф��Oó��U+�B�����<��j� �S�J��t�0�}�������iѧ�pm�;y�i%a�8'[Z��x��w��Ly�l�N�O��@�ԩ�0�K�#=�VD|C�ws�O�ܥ9tL��9�O+X� �ʐ9hʋM�8m�A�L�~J�^�O��W�Щm�*��gw�tћC���.��"W�f�Ǣ7����W�/��H���ra��**��3�T�q��v�o2r�N@�觻v	�-(퀢����8��H!��䡧�=?ǢcL��cV_��Ĺ�!����Ҏbp�-/�K��/�,y?y��:Qd1�w�eS����F�>����=FF"u<(g�G˝7��������v���͠s��e�6ek2�AS�Z�,y�O�6j+��H����H���I�f�фZq<�!�d�������-u��;+��y�)J�ۦUL����eqW�v�/{ÌZ�Z��W��t\Qˀh]���*q���]Z�et���=�N�r&���=�rj>�E������:�Q��-�~%X�bz(��*�\$)�~��k����`�U��b|��'o/�P���QMp�Ȳ�?��D����$k����!� �i�3X#DX�@%�_�Y�8rnq'a0n�D2�5�*
�H�R<�	�a�G���[�!)��� ��?-ȇp�dJ{w1b��mE=T��� ���D�-3��n?��/�uN��.��sCP��y��Y��o=�{6B��E���MJle���E�<�q�j=j��i	�&#�Ѥ�I!t����V����F�6�f �g��W��P�[l^�y�Dh!D�TZ�L���) �C��E;~G�#��ϓﶖ�"{�gxE9���O� ��g�a�P�E�HO?fO#K6����)	,k|B���W��m�%m��՝���M������-�>�������O`�:r�hG�Ty��j�}�A������肸;/�t�S� (ZՅ�*���bF>��:0��a�5O��m��Ss������_�×����l<��� "�ƨJ�`��vJf�X�LJs4.��=�zcͥs��#b~xZ�0��B0��ث��N�������R�?�����I� x��8�!�[�/�\!�B,]QFy��uH¿i�88�v�o�/�4ѺS=eJJ�V�WUGOq�߰�Ј[�&N?��6�%#�6�$�&;�{��x��aM�vK{D��Np�Cj���j����^���˗;���5���!���_���<�T��;l���-�%�c�d+ z�W'� �E��6 N�/nn_�z�Vi�á��]Hsw"���υX�NSi��|$,���x ���H@�_Sďv �'7Rpxq�ו�|��X,S,@��<���!k`{A7j
� )��#'cV	[F��� >�(��P�d>!)�egw�"�}n��s1D{qB�H ��Ᾱky��Z)�J�(g��>Io�_*D��l.9�d)���Cղԓx����3I��4��w1����-��Ga�d����@�#?�_P��0(13��DI�+b�~�G!h��c5�:L��;@~�mVp>|?���l���.�?� }�0\I�F�L��&��,�N�����7߭6+ɕ+��#�'pϢ�	��X��D����L@�
�:��Ōȧ��(�N�B�[��e�3b���]��/u�S�ƲL���#r�����W|K.&�L~���x�H�����H����H��n�������"��H`M#R����-]���`�+�)���5�e��'����ɉS�|�[؁���V=��ʇ�6d(���uW�0����������z�h}h�r}tnW�E|�_��i-	�f&&<�ܻá�#�j2 >w�)�,w{��٣�w����Έ���^R��C�Bѣ��Z��/�������������>�z�����?P�����Gl��\��,
4 �����F=��5GBP��Ae����ࢢ&_�~���
� H����F� \Uǧb��|AHw��>�TR��Cԗ���aw�|��[��!�~��4{�BU@Hm	�1�ze5y���'G|�y�J�i報�)yt=D��"����o��W�~|��_�4H�!>���t�����V�3�^3G`��L9��W�Ԅ���^ΐ�Ks#�A#�\H�4ԏO��f"�5�ͨغ+8��Zӏ�%t�z_"s�&=���[�UKw�����⃊6���tI��G��:BM/(Dl����f��I����1�;�wu��q��L�{?��8*��Xe�5'���!���`l���_W��.����*1��2l�Me�	�)�"e��ˎ)i.�O��8�+�-p9�:��X bQW�([�e8a�4���V�d��Ӽ7�롩�=Q�/��o�z�oph�N7�CQ�~c�=T�q��v¤�%���@Q!Ϭ��D�8l����j8��ӛ���0ԭ>U��.-�|һ�%�-P|��X�x@y@]�@Q1d�&E�$��!.�S��Sņ�Iw��L�y���5�T�<��x���8ڐ0�<�Q�U�+�'��B���E_?#Ŕz]��� f���I��Ó�J&'�/�k]�9ur$�k�,vIV6�A�g%-5\����T�_׉~���Q�ٚZ����n�������
z�>�z�Qa���Z`�Ipk!zb]�,�i9N�r#%>nՎH]_|���Vևژ ͯ�N�L��4�77ւhf+i/�B~��[If�|���S�k3Hv�l��a:"���:O���3�4?~s;��T�jo�7���,Yn���fO���f;-��M��PU*u��k!�`f�o��`Kt�R8=]��U���kL� �t~0{��v��~�P�l`�jca����8H������`���=/�T�@����0�C.r���ӀX	��q`c}�	1��rd�VWcfG��jk�Y��r���Z�f�we��O�!�E����4�&Yb��=�M�4L"e���a�e/�v�I��;6M5��������,�k7}�� �*�pok7-��*,B��o����"��{(�$�Z/�R�A�R�P|�9�6����3P���/�r��R�΍1�ufXs���k����슅{��v�*�J����i	e�*�`��tH��TgX=�p�r���e���FbX�U]�`=3�&pxq{��PτiN�B_��ؒ`�E"o� +���o��ѓK���:v��Hf�/\3�O��IÓt$9�ϐ
.�r��<���0��7,��#._�|e9�$�%��� X+4�֧A����^��7�m�@׬��]^�7�YD�����~�)9���t��v9�"rjU�3� �]�{,��q˭��+�$M����|�H�(KmU'�`�}�����I�Uw���ڌ�8� �d���m��%j��B܈���;���^� V?l_�8�"���̶e���Y������N���}$��?��i��e�)ϣ%�}�m!�%���>�H�;�R�n�T��T4�x���w}%�o5�ʳ�|�=�'8��/��+'�+ǀZ|��%��ҟ�Gb>��鑓����ȏ/���j��V�����g	/��8t��߅/ƶ�Կs�o>N��Ȋ�ꛔ���s�����
P�S'��l�3�6�hO5��VB�BCf'T
5�tD�Lh���m� �|*�_3�놖� U\	6�+�������;F���f�)�B> ��Ҝ�$b�M�C�4�UXa@-�~�t�l����w�J�����ů'���%��I�y
�#t��-�VnJX[��J�x{Lο�����l|o���^����Y:����H�}�7�-��r�}�WAٓӜV�j0'%{�w���q<��	��w48VX�y#}�x��O&������I�D(� G:s��'�6V�����%�d��J_xH��� *hKcs�D�%Z�[y�&P^�<y�"jC�A�o��v1��,��kb�(��?|�j�k}
L RG�^r��a���VLC*g�*loȵ��?8���_�Awd����z�㥔R�aaoQLS��No�5�֯&���KJ��h$��;�]Q�p	z��:���fҷuZ�ժ�dE.!�)�E�-&/|:%Q3/9����'�ߥ̀��H�e;�Ң���?���/�G31$m܂HUnU�D�(U�����ԅ.|+��b�I;��v�>wO�5�< ���B�O��Ya&]Tr\�'��9����Ŝ"�[���y`Dg���V�MDv�2�
Ȳ�aW��rE~s�G����[�RC�e���|�(�įU��5�M���a]n�g�L[ٿ-3�jP�S&]�k�墬�	�¶`Aal�Cz]�}`�x\؉b�B;�ob�-�#hAH�ׅ}����j�@H��>~��=�+��`��%d���A$�Kb���uG�����+��N����d�ƲGU��d[ A1P49���5��l�rׇ�L��"`1�B	��h�@�q4�~c�J�7��0ԚV;ܴ|����K*�lh8&�\䯝�T[V�'�`ɨ2�l��XlxV64EB    9a8d    19a0��TMl�x���*�H�Ƹ��̜�|��_���[m�~"T������K�K�6���u]�
{���#��ϭH;b�$k�����? �Сp�������&�<[������ۦČ������;h�%	y״[�����M���R��N�d��b�� ӣ�$!4�W�}ݙ嗫R�O�"���	�]��,���z��NLR�������$F=Q�p�M�sx�)P.-4m+��W@ivFb��x�;����[o�)	I��^��1�e�Em/&�Z�z�=tn*��%�mze�-m7��Znp�u0���?���Ћ�8�بn�h���n�(����~M�$F�#��5�w�#��g8��.S&�Vh{$ahv�bۥ��n�w8�?��	�G�<�����JF��wH��ጫ����]4P{,?I��X�/Ӊ{%?���A��o+q��dGcʤ
�))����ƀ��!�7x�R��ȣ�F�e 1��P��pB���(���ޭ�Ҩ�!�F]����N4����$���	���enCS��A����e�lB�#�z�H1��V�mF}�U��8��K���`(�/UD����T��YքC�[�\:I�9Bz���
�*ç��k��C��S�kg�v��t��݆St�Hv&�:�-n���y�U����H51�����j��82 �ѽl�I7CޥCf;#A��ͮ��'}�+���{�ܧ���)c�	BQ��*� y�z  ��D�Ji:�婟Q�Sh`o�I	�As�A�b�H���GPR�c!g�P�x4eZe�{s� Ɇ	�\ﻬ���cFy4L[XC��k�:���YPM���?�&e���0[xC�p�,}A�� E��0@�#�l����e�O�[��E�C���WdE01��~�Q���SٰmϬOQ�]$���Tt�Zz�����]�U$?��T�J���KNz!Ae׾�y��б�P��$y8�t��:�-���F��^�¼����
��f6ڷR�����v��n�ҞT����*bN���=��,�G�Ӄ��T�����hܬiv�z#��OL;��^��SD�>�R�J��G=�7�2��)�.�_�뾉�I_���:���T��N�Y�/��J�>�z�B9̅z��g���8�H��$�����U�gM�r~���qKlA쫔g-O{ ��ܣx�s�z�j�v�f��B��i��t�$B�dW�o��5(�,�g���YӉ��ޚV �P�=T�fm���+�1\;����`�Qp�֩����s���e�d�yh���EJ��\�ł���#�d��P��kk�l�33���}+�����7����8"D	�b��퐜[P�!�����H�a#���gTAd�b�^`U� !�=���X<A��Q���f<wyK�C��ֱ\���IACۮI�k�<UA ���uE
���.'��oҕ�@LU�@Z��W7�1޻:*m\i	˂]�%qE����az��`���]�%X�n���ǻӪ]����� n��Z�.bCrhQ5��a�m�������u�Y�Oy��Y�hӢg�n;��j����2�<��p��|�V��Cj* ���Ok�������t ���R�t��D����� �.��o�@6��}��"7�t ?�b�����̻$���yj@qxo�
�WJ��$YRn'��u�;Yl@P�s��K�� m���}�D$�$q��==�[����M�w�?��o`C��^]B����"ywS�5�w>sm�����W4n���{w�JSgq��^X��l�4y�-��W����n��/�);/@l�E�J@"
/�aq�����sƯ��QҠ�<JS9I�YV�up�� >��DGF���B5�q�t�J�ޜ��� �)��f��M �?nG.q�$f6�3��(|��h���D�{)���OS~W�F,��ԡ�I��)�?7���@!�e{�H;�)�l���%Ch���l�������p�6��w����Qװ()D� ��Y���N6���	{#v�OW�/ݱ�E����ҙh�����?	B�Ӓ�����9�~#[:J�A���ͅ�8�)_b?�!U�|?�ӕ��.�v�'�_t"��U쌻�z�e�E�d�g�A�~��h��0�S����ϧfҀ�����߁��[������N�����v~P-L��C�����x��#K�"{�]����J��.#�0�����ƥ$�l���j��2���70i����Cn2�qA]�v���y�\��^���FؑO{qu�[_�*��C ��NPg�]����"������D�A������Y�煲�q,��ӧ�xsߊ�������>prP׮���1�ߏ�93�Pͮ�{쥺�����i�OMX��G�VK2o�e{|=Km��:r�CI{�s�6e��=�B�)�dt"z"h��\�1�/�V&���Z�#��i'ʐ�q{�y]�H�=�׸Oߕ�s'� �K���jd ��s�@�-��(�j�M���+4��J�����i6p��s���c"�&*:��%ґ���0S�;���-�\�,Y�o4�:��l���Y����i��s�%�~��S�%�3����aƟc�����#O�Q�ao�6-����>mY��+�s��G��(�^ǘ��\4,����O�E�b�L�l>��n��MM�@g �}����Ȇ�;�k� ȩ��]��0�G��+%�7f����dw�.���NL��}��
����w�5%���絧����$_n�ڍ��}X��]�150���Šx�����=-��NC���nW��=V#�=De��W���\� ��Ki:���-�_��"��y���d%�t���+�X�;��jL�ñQ��Ů�?�9��A��¹^�5/qśThك
�8�nG3��:�}�|�P��C�Ҁ]9��ѯx��y�ڦ"o6��>C9����:��*_��/jj�	�a��2�%��כ6����d��Й�����V�K��.^��)�5�Ka��7��E�w@�x�T��6ت_e{��G���|o� ;#[c?�� ���R5�=���ٮ�eK�f�8Z�B^�(8m�����){���Ē�l �W�>���_2s�~�qЎL.�L�`��q^�bc�-Ԫ�ݯ��A	�DW�����o�Sº��0�u�	L�;aw�,Y�Y>{�h�4����8��d�L�v���n��e�没�;����H�UқG�� G&�E^1��[���%�wXӛƭ�]\��Z4���h�x�\?�@ꔛ�����J��KFH�]��L\f_�ĕ��)$�5s�z��	z\I�̐�h� WLX�7�I�d��Yv����۞�$��LE�w��.8i)����f���2��gg�p�8�x�:G#s��t�/q咖D�2�A�N����M�h.l�Z���n�£��y�u��c=xy�ǃ6���5�/	�tEX��ܬ�������z*������]~w&8-�k/�'&J�ŷJ��6�W���kM�=xb�7���[����#�-����mm�Uq8Z� K��ps��#Xv&EEU97]P�\���X(�l�d���5\`AsP؍��y�\|{Lb3�d7����L�s
�ԙ͓�ԫ���v��qr�2X��f[#��y���/�Q��u��\�D�(oi4��0��]�_��j�'�X��INҟ���e}뇽I�Eo�Кe
ǆ��uf#�?͂�䁀�Ez�@�ҩ+u��=0[�{��P^A�*N�5�dD�r3=�06�c����q^P1!������vG�T���颧jxa��b"����^M��R��5ZV�:�&¾c��u�h��L~
���ص>y�F������U&����Q�#-��E���y�2X��� hN��|��U��bV��������L��o%'nG?8R"�s���&�U�H�7� �	�(�]�>0P�o�-}��׻�Ars!T	��� 9��7L�Ķ_���'{�[M���W�����8$���zk�5���v �z �<��
:wbf���o���xh/E9�}��17� �^en��؝���HW4���3]�yٸpi�?�"D*3�)��]w-�	OE$�9�O]��y��5 ���Uxu�Ib��˲��_�V�r��&��#A���Cv��f������Y,��%�ڀ톲�5�y��k:����b��$3�� !�O6�����kS��H����:��S}����D)}a�K���<Ԅ ��"���śM�i1�}��t�]ש��VE����N�Ы�n��bݡ��0�f����[�@M�)5�x�9z=��~I�r�m�7"H�^��Y����L+�k���.�Y��J���j����Y�G����#�j6����mBs�߈�6+�N���S����Kζe�O;7��A���⧑ZD(�eC��0GTvb)�lp���'��8�,�8����nߍ�p�8�Pl�J���D��F��P*�S��Y�x@��D�t�É�,Ls���!�ij�꧜�b�1�<�=����3Kޖ�����~C�@ؖZ��}Y�Utx@����q�j߮b>�f��Q�&EF��p�fu�L�/�+����bA� �KCbeoo�E�3����ŏ�������VC�eT�G1&L�t�s�ab�k�fjE��!�b{�D�]�l�q��"s��M����>�.�ͅ����5r<�4�#���#��;�n�4!������^`Bl�̃�JbD!6��X�~ �r.��']7�/lr��#��)ɨ�(4�V�q��?���hm�x��(X�u^�+��K'����T+�+�>Q��D�e�R߄����[p3co�"�]��"у�*E�\�=� Vݾlxth�^޻YL&��=k��Xn��&�a -����A���a�'�Y��	���kq�S�eN�ϟ�v� M.<���(�w��E�"�w��j2uA�g�I�mѐ'郖w��G�������S���XC �a>��lV^ka���;�k�k̬~\�VDA�h��Q�뜽+��;+Ǯ�޴��eq�S\��0A�R�����e��q��w�`��@���S6���&2'f(���x��N��L�=�;�"	&���k,sv-���.��%[���ҺX�$ �	�EΖ˾D�2*[me�2�1��.C�΅���T���x�� �F���P�f��2P�V�2W��|��"��� Û�8��=�b�"�,�"\|��)�ujk��q����
��(�I]Q���@��z����J�8鬂��#����W|��2p^�*Ȍ��k�h��lnv����64JX�^)�q%�.К�qI�[�����,�Ԩզ�5؃���{Um��sF�_�����r�c��m��u`O�"y�i�y
F(,�����WY������O���z��~?����ܕ/�U���*㨩���y.U킠
y g�����ǻ��_J�gɓ����[(1o�(�)�o_�g�;���t�5Eӌ~�V"�A8��!���80��Lא�-����T���uG1n/���<�R{����ed/Ϗ��� %.�&���;��x�'��E�b�5��� �#��b��s�;���
��S�8�[��A����J�fs�|�J�U���������
���ߋ� ��fہN6��c/ox)��1���3�ר>��ֿW����ܙ�EŌ[h��3�i�)�j�'�-Z&%��ʹ��ۚ��:��K��+c"��� �j������8�R��(7$~�@J�а����DBe�C��6���n���_�S�l��y �؁�@��n3����F	�Ԥ��-�O/vq�K��#W�ǋag�(<����ւ����]F�`��B+��R�£f��p=g4Y15�F1��%%���}a�i��z���ڤ������T��Q��͂�?r-��:~r��x�T��4Q�1�Ox+��=�z)y��7��V
�������� @,�m�������~�Y&�ILAb6�m ;#�&yHC�4�X�z�C�w�|��kSq�[)�&����kmD媔�!B��o,��F�p�b%W�J?�y�
����+�{E�� E%D�y��|��Yv���m��8$r ��K��eQ*���`� �$d��h}�PL/�f��ۇ�s�l����V��s�����DE�M� 3DyP+�9{�����>�R������l��C���kH�r��fW}{G�!ʒ���#�W��#�5�ea�@����]̳��5���A�a͟�*�<ٵ�lp۷�Z|{���MpS9��\���<�Ȑ3�#� _7��UB��R�Lx�^��L�a���9�xs��"�F��l��]л/@.��D������O-&N
ũ:�3.g����y��4�`�xA�ms������c�����o��0E\�