XlxV64EB    20d7     b30k�s��̸I6��M|��C�ξ������N�*��G�#�AD�V�\�uA�������ل��B������?)�D���w�����4�^I7<�R#K��ccYp6�����qO���-]��e�'�&��r�Z��VpD1�؆Ԛl9�$0���+ 9[���
��9��%b�� ^ZT�ߛs㑓V�X�+^g�wN�8����i�(�k@��l�������*���!�TcOm>�Y���8'$��:��>�pL 8d��*�n}�����q��g�\�0�8���u��E�B�����~�ށ
�R2�r��ݶM<�ޙMV����)��]>�`z���t����`�P�vT����K���N6¤^����}#(��(/���g$�!��U���茣C��n�����F�����8[������Ⱏ`+X�g$=�޷^A<gl��dhՁ�� �p股Ϙ����顬��3@�0`��V\J����,�����)��]�o�1����ñp@۾��B:�.��))�0�x0��K��J�U��+P�Y
5ʰc�7��r|�)�+L��V�c���#|fS]dz��S���S��Sf�^�w]�����H�L�I:gP��o#�B7()��
�J����{�l���:u�����w��(s� L-m.�Ċ���֋L�5�	"
�`q�-� B+�r�楑�OnC*;14��[{X��.rn9���q�y7H���0f�h����Vީׄ�?���!ʹ�J^�n��+"���=0�.��0#/So��p�P���T4�c)`��Q#Y�O �f�T���鷥�:A#U�^_zf�Œv����
(V��v�+�}�I�>�F���<��'�~�@�����.O�]��z����B�&�v�Ѭ�������Z��x9$U���*���;k���)���l5
��&��Gֺƞ6�,\+.����"V1n%�\[5Xz��m,qf�
�£t���$��rj|���x�Si�슷���K��	���⾮.ڄ��Ms�<��Jd���Zf��k�/㵺�Zq�x��ZZ�έVu�K͂�v`���=�\[bz�XO�&�cg��"���ӫ��d�'�~؇���b7�����|��6� �rT�UV*ϩ;�\1쬈Q�zttp����!Z�ǣ�S�v��$����Ro~!��^�䈦�!��sX�Z�6�&W�yqΛ����txW�D4~l���ݔ�"���l�n�F�7�~Tc4��U2/��^�.%)��Z�eI�yV@�K@	�̊xG�l���N&�𻁶��P%w5'���%J�0gr�	��j�̸� LaM�`��s�4��6���{Nq�����ۙq����O��+��l0��s�3�)gS�Gf�p_��zC`���������Jψ��)��V��?�?;n>vBib���b���
iA��P`�m�[�Jh�2�c����=͙^#�.oC� tJ������JO5���;�V\{N�q������Ze �ɒ����
ɢ�7��Ku��h��v�k󮭝:��>�ka������	cc��'�qW�q`̒w8���1j�����֪/�>d�Ή� د��"�a~��D��[�A{S��`��6;'�Fh��QD�x�m��]�@�M��m�Y/x����*���'$�:6pƒ���%���<���� U6�KH6Z�A�媼��H��\�z<כ����]#��o�^<�>��-H䗅 !�x�pã�Q_(C��J��;���Y�EU�XRT"2�}y[ �"��Q݋���C%�Q�ف2�����?Z/+4PVȷw��Ѻ�s�\��B��;��ȭe,�IX���k��?M���܋zqjVl+�\$����8j��H�/F6-����^lB�=�����#������:��N�c��)�}˴I��1��Fp�#؈��˜QOr}�\�i2�tA�����!�k�IU|b�7���^��?���E"Zw�c�u�Պ錖�a��t.��<vJ��F�@�{]��O��:����Np�Wg�N�-L 21�ܤ�e�F��?J-*c�cǭ;��L�}���f����xl(AEYh�:B)�_`�G�Pu\�U�;t�(�����yk�#�6�2@^?ࡳUleu4���w�E�m���Jex1��	&����	��5v�}Hb�vI���5�S�v ���N7Vt%}��x�p�Xi��K��\�U��a+do�)[����V1Ztc�s#Q2[SG���JN��ѽ�� �U��f쥛�Fױ�Pv/Z��"��'K?��A@�G?��Rc.�	�ϛ�^���A�)v�'e蹠s=8�"H�ZW/���X��h���Ofp	���z�-��%�-&����f~'�'U%	$:�}���'U;z�=�ݜ�הí��ńP70�&T�`%�4et��b�IҦ��h�L|-٫��ЅC��*}+p-��p9dh����V|������½�[K,ˡ��DG� [_��D���)��t]xȞ�t��_�TR��*�hH��i"(���}�6�d�����7Q�>��5[qL�M����;R�����˾ô��_'������g鳉�u������>ȾU�/����~����Va��yQ��6|B�!�;,b��{��k"���1 k8.2��>Jad� ��V.� ���X�<��2)��y�b~hV�����1���!Ω����T��2�Zʃk)9���{��w��ձh�m�!��M�؃h�	��:��F��I؍f��Y��A���pӆ:�����=�!�p{	p�;	���Gj{,&�訐��6o~