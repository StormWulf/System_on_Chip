XlxV64EB    517b    1220�*�����G��*�Ш�}wV�Ҩ��L��l���:>N��d)��j�i�O5u5�'��5��aR��:"�Bm�Sf<}��e:��	��+�Y�Qx��� �n��9�
![�����Ўv���B�T�ʺy��4�ʔ��E��L�,)�v�z|�� ���w��]��:bo��+�&�E���#;R�<�	vPe_�+����
[;�p�M1�H�n��a.JK`z0���ᛢsщ��1�
r�}���$(d�,N�Hqp<��H�Ĉk��fVq򪧯��t`[�1����4��i�����8�CL���o�g�l
cs4����6�z}F����.��(�3�tP��^�2���bB��D!s�����q�	��o�Aſ	��.��n�KW��9O��A�T{��h�,t�J�N�fJ
*[&I�kر}��ܮY�ަ����y ��Z�a����O-I���ݯ�:�6/���ia�3Y�U�U�LW���� ���Dh0N����UFEFO�6Ox���e+z'tR��k�D�����j�M9�(l� ���1�㘃��̐�W���]�X͂��z�E1םЄ��|W��f֔&�kH�]���cU�(.$4It֐�d-��e��m�fR�4[}b�`g��d��=����[�{�P+��W���5)��	R�u)�:f9����e�f�"�����]��7�u���U�x'��C��,���0W�Ehv��sNx��7�9���:\����M� �כ�_$�^�<F����*��y�m�]���E$*�i=��d;[H⨴I�r�6m(SO�L�ST�����	�3C�ߨ���ׯQ���O���H�?:��d��X�"۴�YKv��߰wX�忤�8«>��a��=���7]�'��>��,"k��'{P���F.�`����x�o=}�.�}B��HIC�H��� ��~�a(��|^�&aq!$=��:X�m�"p� ^O6v/L�;��o�����ܼ�=�����)��F���iN�$�ʽ`u�'e3�rkX�A&0F,���7lP�����3��vqj���>�R	.R��Ka�l;z�'���n��j�<7��j͘L�̫{J�bv;)��`�)���(��^d ��-��!�-���Y��w����}�ƒI��`�����s?�3�(��r�<%��_�\����QƛBN)�Ie~�6�6�0��w;��*L�s _�����|R����"'�x�m�U��]��ǜ�\���x<&��o@ZZ^�hnR7`$��?6��C�U)��?�i�L��2�L]�Q�'e�]ܰ^.�%i�1�o-Uc{�Cy��x�
��W���:%߻���5�-n%c�wQoG���t�������yo�]���_U�ּZ�u��Fg�F��q���UɤPq�iCRNR��O���9n)}N���s�R2GK x����1m2�ױU=���N�Gj�}1�w)��-J��m4��]�>���^�]�'d
�#ǣ�}N0�ˮ^G���a�h��ȍ?w��c=�膛5��k�$�M�v�qK
�G��׶	e�N�UQG�;�0U7�"��#�����1�»Fy됁(+�U?�k���ԥ�#����J��WMc��K��I���E��{��J��_p,���0�b��oRzs�q��^q޳0����q(v�[h��I1�`S�x�7L	�	W�n��n���j�����o�"��,l<ĸ��~j��Q�@���g�J��w�4����h�O(SA�(��{<ǩ5#~�"�\��
�Lk�ir�H�q�X�*�<B�`��Ey5��U�JJ$_�\_�QL3\	��e�o�i�"i��:eU�r�C��*]���0�"�GҢ��9Bظ~���p�ܠ��ոպ�計�*������_Q�df�l��Z5�_�����k|���x����l�H�="c!�s�G՟��מo��?�mt����Q��)�
=���:��-�ũ�*k�4׍��\2�3.t�z �X��ꅌb��6Ri��16w�_�:h�n7�u�g�l�f���W�@��z̓��Z�LR��=j��g�%�L���|λc	��=�gK��D��֋�q��H�E!)�O�V�)�QS��x�w硍�p�29@�-c�@���H��y'��-�"$|���>�s�9<_��.,��R��͐.\�E�x�u�Gl�8-���O�;��������_����X�ݩ��1A��B�t�m�����U�͘���#�K�;b�,�͆+��+�%��,��9�3�[~��o2�<����9�ኩpP�Rnv��dv��_���L�{���%�G�Z"w��,���4�q=�dN�) 3
�G�TR���ԏ�#Z�Z�<(�s���ڈ��|V�>�L����5E�Բ�ROE\�c?ʣ�pT����Y�Kn\Ԝ��Kv�Hm �4䔽���3M������؀^p�z��]窶4�.���gm�k�T:
���S����ԓﷁ(󷰄�b<K�!P��b�pݗ^��$R�4��+�7����B*��ě���{(�R��R�j���3�����0�ȱ`�l��u���S�L��}}6�k\"�i��Ќi�+�c�
�a�B�_�E�/��A}��RW^`H	 ��R`�������%.;r�Ȃ�-��Г�Ǒ��4�.�賧�l�.��&��f��^ִ���.ǃC�l���I����a��D��!��	'��C�ۂ��ۓ�t��3��1�P�'+^^��� �����L�`3Von��|X�(�ϏK\:w�[6`H�k 	�����#��(Z=ALy���>X�����<>��BQpΚ�5��8���YҚCE��?�_���I�5�KoZ�,*�J�on�����3��R�=6��_��T*5兣D��t*Z#g��M�J�jጤ�C���X�ʅ82��U�i��7yG�,i_$5�G �՗�SbVh �yȅ��3�r*�I7p�HX����o���a}��i�j#�Wo�P�R�w䛢X����j~j|y�=nÐ�]͍��ۋ�S�2���zԡ>:��(̛��0��[��Z~ZH~>� ɬ�(�".^����"3�Y�vZAaW��ǚ���0Z�����<n���u'��Dp5�Z�G��wd�5 ��J.��tF6Y۝�zQ�	�{���T�Ӳ���8��x���Z'  ���`�LF�3ؖf���VcR��\j&Z�!m2o)�"�u��}��=ڟ_+�Κ8��n��0i�=�Eo7l��hSd��}��C�3�w���s��z��Ŕ����pr*�$ˆ����W��S0H�r�aI�����krx*ը+�w�;���zlI��&��M0.z���ʪ%�E�L��M�R�UEy�l�!�ژ���N�_�z�W��DLOjTd���!2?=J��t[��D���3�
�-<�zׂL��|�G��C.b۹[�`J��E�K�7%�J��;&P��y��=D��M؈
Mi?2^����e�� �=���1ƿii�_�z���O�K�2:�������8^���*�@\��x��e��0��E�����Fy��y��}ʇm���M�*����d�f�5)<\�*7=�A{1�2��Ä�ł�2+2k	�\@wR�h�oU��]�q�K7j�	m�f@��J��U=�2l�$�Ͱt̽4d�#�}�+��y/5vܭ���z�=�L6D�n(�l��A�[�R���Kf\t�lE���$��v���$���]���-�p��B�*YOo~Kkױ@�+0��?0��Ԗ���qv�}���5#`]�c�W��ڽ�ri���O4h*'
�s��TRuX��|~�j�C������ؙ���g���� �����_��r\�60�qޝ�;{���=y�p�=6�㕥&��$H��?�a�R�r�/���Zu�`���%����@�9�!�:'����0�a�G���߷ط9��4}E�܈���+ss7�PV�|�����������>��^ʹ��3lm���
H�s��Gw|a�.��!ة�Y��}> �X�jrtc�;_VS;_l�x��\%}M�d�xl���ڈ�}ʅn���it��U&��ݘ���a�j�"˗�LD2 $�f�R{����2M9h��ͤat��� ��I��1�5�@4��8�
��lJ��*0�����ս��r�;���9���9BYG;�:Œ2	Pf§�x,�TW����<���sP5^�g�d�
��jSu��
��������"1�z�06s,k�4�H*J���]r��~�,��u	�&b1�3Z�.��������Ds��,�b�ֳ9����]�$F�W�i��&W7�R<��Kj�.c��2� 0]>�J<29�u��P�^0t��p��Ʉ���Z�Чcb꠷�L~�"�n5�n���Û�,�S�� U(��ݸv>W�t�o[O�#+g�,�6	�
����m��([��C������hk~џ���+�h
Te���AJ��ī��,s�j�/��E��-_�]��&=ğփ��������>?b��TxL���n2T��