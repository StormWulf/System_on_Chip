XlxV64EB    1681     8a0�r��q��>�E�bW����@�t#TP(p�,{����Z?Tx~+ 0�ӰXtZ8,����d)��Vf�i@�r��eđ��Y��bm�N�ӷ��T��q���oR5�f-������>!�*i�a4��nց�[��|-)ŉ���x��6_>Q�����Z@י�3���/����kT��*���"�£īp\�i���}=ݢ2l{����CV�lo���<��'w�&Kz���g�0%!�J�����>T`�\��ew�,��a��8���5=��!�Gc)���[����&��$� s���C�"��.����0<�,�sC)\!��ϥ竗C��w��)d�+�ܒ���́R�T6U��ǮY��,vi�x�x5e�O���7c��E��}��\$0'���^oD=�bי�i��\r}I�e��3+	��uԖ�u*�WB����r�҅�w�����e���9�Jv댚���23��s�NJ�WLG�6��)#�M$��Oٹ�a���i!�S���Ҍ���cd�N��A8����ekoa=
Zwp"uR� 5 *��:i�F愯P�F�3wW�0�L���G^�:܊�]�ţ�������{��}��$�^��-�?��u�{��$yWY��8#��Om��VE�c�D��~ws�QIE��l��MYo<*��xE·�8��(�ۀ{��� v��uk�
����o�:M��R�w�@��� Fd$@g�����:y����yp��Bx�-�����vt��u��oA�cŭ�R�g-��*z��q�M/�}�}�sR)�潪�.��!�S
(�d�ξ��%��s.�q**�M�}�#���O���C��R�M(�h��F��g�e�Kg@#h
q)�1~��w�}1H4�s8W��O[K��0�ߡ���)���'����W���!�SJv�Wx#���/� �*(�������4�_�.�O�3�HM�d y%&.���9/mG�4� ρ�Ӟ�ol�poJgs2פ��^�� ��U�ܑ����k�2�AضehC^���}�1x	��r��=}y'�
�km���1"���O�`Hf4����x�0=�})>6��A/�%�k�$��s�2�a	�21��3��������h����GY�:��MM=T��F+�7�ݏ��q.p�H�e���I}����zv��c�����4΢q �4�u b��}���W��i�bh`����w)�1�������]I�:��Ƨ5٠��d���|Z�-�ׇ˦k�b�cE��)�d��<y��b��S!y��5بx2�˶���(�1�H���kQ�������'F��k1�DV��<�;;K�8�!_n@��T��R�vi���!'�}�>�;Yup%bV2Y�V���j��ʩ�ea��+���m�9����v��
��x�9��iyK.��F�y%b��R��+�3~�NyǮC���e�V��t4��y�m'��Q�wK�?���9u��������l�h���%-Lô#f}��.�%�|F�4���B���(f����������曘˕V'�c��q���¦�,���2���yP�w�p�1x�B�;3��u^�~j�������#~�R1�$��d��7�K��,b{�~�9v��1;�J#J���?ɂ�vݧ�1jW�r������7U|����ہ��Gas	�lsB��	ԅ���;&*��C�B$��$�Z�Y���:�x�c0��<��?�r�%�JA"K�w�i�!����L����r���Ȁ�)f]�:�}j��UA��ڔ�d@nZ�C/ha��:��'���Q���1X0�F�L�m\s�|�:.���� F�#,��W�Y��?�F�k������$��A{E.뚱�!D;�̿��
��/hܹ,Q�[��k�裸mĠw3���B���n�*qgo@ЦV��U=nA�ӂ�9��t���V򊨋��!Fa,�������i1�m��i:�T������Cg���_��$��vǡM�t}�$�y�D�g����j��t#�s㐭X���4[��%`�	�ҡ���DX�]�u)��َh��l;��`����(�t���j6���أ�D8F��|�6J�!Q�u{�N2�E�r	��.Еe���{��@h�;�����a���v[rf�iR���i