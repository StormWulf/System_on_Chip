XlxV64EB    fa00    24806\��qY�,IĮ"�� Z��9��4 a�z�?�Q��?���?m&4�� ?T���k�Db�o�'�ԓ�ł�V5��\�������&�;���e�Γ�7h�� �y�A��Ca��EƩ���7�=DO���7�(JpI��k_��j�D�h�����T���uX�u��aF�,�JI��9�+�z.o�)W0N���p���Π���&���޵Z�^P�j��+n�]F�h���k��P���ͅN�.�����#�m��]3��V���>+�U����	��Q_
�i^�&�"z�T<�OZ�6��yv�0-����,^&`�2Q鵢ܹ��BAR#����T�M&M�s���}4�Ww�D���5���x�f�^��9 ���a��6{���{ve.l,�Y3�x���ص�u#95���k�~���LC�
�-��5�hzJ­��IuT���n_-��	������w�u�qૈQZ�SW��彳�I����Ȏ�C<`��ɓ�m��=_��w�ָ���ϱv��2K�^�R؋�\�u��0c*�Ծ5�|�ٵ��	LB0�%V�W,����`��:�k�JO�G�=�,P�H��;�翠�>��[�@�{xK��)hH�Iw��i� ���Z��;<!{��Bh�G��7-uB�~Vj�;:V��$K����8N���iV�x�[���R)�����j=�
�^� �ɒ�#�%�q�g�b����{����Y��s�p��U�My)��GD��׃Ljxc+�ՙ����Ƈےd3.W�^�h/�^��+=0�\x6YTéL���VO2�]�BɓzN�c�BK�>����	�c��v�����`��{��o��M�i������V����h�8��㒟���,(�l��.��6��&c1�x��i��a��+)M,��L�B�KeZ�l8�v��\ �B$�����i��L���h��P~ب�/�>)�k{a������vqS2vng?��*Ca���n�-���L�g�5*X�`a��e���b�t�!�z��f���s�D��λWR��W�+�����+?#����c��ؗ���|����I�Eد����Xq`6{���: �)q�<�q�[3Y$�"d�*xU�֓�	�#+\�ԝ���CF��������u�������-չxR�Fg�⻣� 6�|�Ϧ!�c*����]!�+}���X��?\��j�9(S['�iH�����RL���
�4>��%����ռ�#!�ꉌvC���ic~��&ᅛU�/�I#��ڷ�I\�}$cb���xh����˚�w������)1C�r�m�aI��~��(�·��8"W{��n79�aS�,uo�X��t����c�xvV������ɷ��Q���t���N��ח7��9\�Y��K��ب����̵&2�-�.�wJ�'Ŵ鄬d�a�}�&1����m�K��U�za�W��SЉ":2�.~��փ\��C���+e�8@��
��$�yf�AI፣��x6�-�#�;�f�5{��T��)hyum�塣��
?���Wꤍ�C����Ӌ)_���J4,0C�y=�LoC4c=���R����g��S#�p���K�?�Mϰ� -v�♊�8b.�UH���T����P�Ͽ�����
��C�/��� ���'�W�@%�U��@�5v ���(uF|@��fmF�U<�����5i�2T����Mhtr��|	񃭂3ҩy�En(&"��5"Δ뷧��U��*H��C���vd��_�8ê?��"k�#05�ЫZ20��ID��.�k�AL ���~���?�v�z�C�ӡwO��TGaQ����UG�I��z���nk�"ϐ:�3�S�,>~�mʬ)/�\�H�V<����N؎���v��;i]H#�4��Y|���L!2Χ5���_1_�+C ��D��qx���K�El��VngÚ��q8��@���%!r|��ҵ���^�-����9΀^MyGb��|�@-*���Xvɚ	�!^�nPt�I�Ja`f']���h`�9;x
�3��]]D�m|%�@Ё���]Pg�
�Ւ���������-
j9^�'��H�5�/~�hE�ԓ�:��"@��I��5�x���ǁ�ߴ>����G[l�	�Ka�5$�S0$P�/�x:q9�� Or� CX݀.���!d#9����Mֈ3BM�����)�;��/u��؍��-�M���ٙ�������	���y�c� [� ���6Q��۪��M)u�������mg��͆P�$Q��V�bal�����WF��$aO�7�`�&���j�
�*q�����;z��v�ՠ��L�6R�֖(�l�e��`$�n�; �p������ sX���o�r~�_���ɶV�V�Y�P�̡S��#�5�'��I��ޘ��n�2���R����r����ic��Ǩ����lx�אw'C�r�"��҃��U�-�V$eg�"��糕TlmK���f�9f�wQ?�fnZf��"��A�j�>=���b"�g�2Y�R|��S�O,� �8�h7߃鼃��²�ؐG�P��NL�*f==�c��n,}��2�=U�l����n��}���n9q�w?q*��U�����YĦ��B`*R(�&I�q��)�?����#-���l�ȥ'z�(�ܚ�t�<�ĭ�F�Y[�50֌�nBX��M޶\�\�$�,�;�q�G,R��˚5�-*���:#��c�P":j�"1=2�@�*P��8�}��IC�v��c�	vͅ
"�m���(���L�sXW� ��y�*���qL��c�x�,B6¡�{�`�&���֧E�/v��p����16�����;�/.�s��n���5#=A�k��Kv(�`O�]�0�gG[m7�� �ڠ���9BIέ��O����8�����߳�) �^���ڒ�* �D<]�1z��=��a�̛s�<#C�٥��@/�V"��c����ܰ�~-���������	�1�T �&��I}��1�]�[,�������T�y��H�
��q˞%P ���xZ��-s��K��� ��q]J�AFSt�N[}�طըx�o,���.H�zZ<�C1i>WTp3�jHѽ��;���Y��i�����ҿ�'�f4M;*�1x|���5h>El��\�f!�.r�0��՚1��T$�h���X0�\j- M�\3�58�t���i�[C��쭐N#Ɠ�#*T��I��ę��dAC1\���Y�$Z-�1C75�Z�*�Z¥ܞ�f����䱰2zOX�rT5�*��%A?`����4#�����=�L�y���ӧk#�S0H����@�K;�Kx-�Y�	VMRz�%4�-�2�Ñ֓K�n��?�YyWj�VΞWi��#��\�� '�%?��
P���9�=p�5�ܗ������m��8�6ZC/�O9Y<Q���j��zl:
6�Ċ�=�S���y:bd�D��b��,*J75Ep�s��}� �_�v�F�ѝ['�����j���|`��}�I!]�5/>�����	�
����-��+�_�V�sm��S�j	�#�S�_�Mjz%��G��O�ET_���U�~A[�3�<7�MH\9�c*�m�X���P���]��C���Df!Ě��_(�e����7{�f$��p����#�e|��o����,�O�R��	�@|�]��y)�� ����旯n(��R��F, ��Yi��\��Q��j���"��N�����m�X����ow�1�����QpSG Y���w��_�;D2꫽VGQb�u�V���2K.bx�T��Sm��Ӟ�*<_���19ʎ-|S��>U�&�գ�O3��V���AijW2��9�?	_$j.�9�Ʌ���C �Q$�,���+�hZ�����R<�����B�s)���Fɋ�"{�����ޯ��W��w#�#˓04�d��wm�b���P�ފ`pS�7��U'ŒU9j�A^��<���4��'1e䋋�͝���������ʙd�r��yf�})�
����7n5��_�M��"'mj~��7�j?���{�����'q�v���0d���ciw+-h��
�c&�N�x��D뵟��r��.>����j6$bޑO��1\��/.������$�y�� I���8YB����1�8���\�����PY�1}�
�v��3H�qf:/q6��J*y�'{=��N�+��
���kL.eKd�vGE�����Hپ����'v(�����?JH�F�L�tD r����U<0��u�׶�~3����ن�Y���Ƃ
�Ore���~���ڈ�B[�d�$Db�"��FIС�CAuaX�b����ܠ��אm��{	U��z�aH��WՓN768KL�������ڣ�.�Pǀ��������`9�����&�SV٣Z�9��Ǥ�U�"*Ȩ��*_��t�5�^)����s�Ѻ��y@��D,WG��N�'U�����tl�!"����\"ͥ��+ƢVs���w��a�� z}g�L�Э�QyQ�qfK�� �V&{���I��g�n�����JW�ؽ���"�f���˥Z��/�?��Վ��Jȋ�����A�f4�	���X�9~L x�z낊Q琮�ˣ�kk}�+;�觷�'�I�y�<������F�,e�,}v���j�d����z����ӼvA�j�uPJ��+��X	�\�N��C����a�R�z$i3�����QY�� ^Q��3�����H^KDio��/�5�y.I^������!{	 �*�$�|��wf���r 0�׏`ZC`-}qH���6����zH�|�;������dr�Lr#|�������)4YwA��lC���Ă[�ֺ�,}l��_]o@I�"��5�� E|�K:�6~���ހͩzÑD8��@Ng�森�Vl#B<�~�|�M�Ǜ����	d�[	�̝�:�/m����&&C����J:E��8#��5f؉�?���#46��@���k?���L�];;Ú�0HQj�֩B�;�ld %R���~q��=*��6�T�Oh~�A���T��_w����\��z����h�������.�Ź���Zo�C13��8t��z$ԡ���0x,�ǖ�;�\a�*`D��h7n�0��M�D%f��_r�s�� h6��!�Ҩ��z�'�dT�򬝹��=֟v��z63�+�Dg�R���v�a�]\/�!N5����_V"j��C"�|�L{dq�Yɾ�B#�_׺?��l��@ �z;Y&����=��5�%��[������9^q톿���D�>��j����������w~�ύB8�F�#�n7�N�܂5�;-8/�|!�~n]�X(��!�n��Η��I��plx�&�0h/v��͠	��u4<iO����GJ��x�C�T ��-��$!� H��Օ�oM0��F���#q��L��Zι����ʎ�ҍ�HmA.'y����5)�z���-��D����R�z�_����!Xr� ?O>�M(u�!��=#K������	Oy1�a�����Fp_���j/7��ZG�+��i�esvIW���m�l�S��v�V(�ߑ,q����df��îĿM�B�ϸ�����	+�Q��c�������@s1��ˠ�������ąǘ�\ev�^�=�{52ӱ�S�HHt�	X�:�u���n�!A����`��k�K�\IuB���Nt��|cе�.��!�I�lB�)��rm��0�Lꬢ���#Dc�>0��/�8�7\�gj�Ue}eE����!�u�䭜4��lq�)�v���VK �1c�ڽE���'�U�{���f�T	�]���Mɱ�Kk�9��7�ҕsMm�A/Bv'���:�(^���E��hht7|�sϸ�0�V�;-y[��[�`-}U+�k9%�� O�&�!�c'���F|����������P��'Ü�P�$V0���.��-�m�nǜ�
ԧ��BE��O��8��e	��E�(�ƅ��xcI_N�R�]�Ĺ�� ������B'���b�e�C:�`��P<��k:n\`�I��A�2P2��x����pyL�wQ�Q�G�gwm�&�3�h�N(����J���J��T����4]G��ت��x����2 t�h���������W6`0J��0|
5ѽ�GM;^����\O��ܒ˛��M�Ń�<�_����k������@�U��2��a@�������Ӈ���T8����}.T��d�@²S�
��d�E]�W�߼t���������uZF?��r�TW��H���1F!�rR��S�S$X���$��D]~E���j9�C�w�o៍p�Qܣ>ޫ GD��ZO��m��>a��t3L8���J�5V~swqȔ�6ah���NF*�oh�V}�k�Մ,� ��+T0^��1$-�;Ƨ`����
l��|�'�o1BV�
��Em8#��,K�V�O�C^�-���5�h����FĨ_&��9CG��ԛN.�&	�^��*�!�f('E�Q��:�="VWϑ���IlA�F�Z�J��ֽ?*�C����4�A���U�
��{�] ���T��t�#sr`��ۣj��� O�M<3��Si�a�{uɈD��Zc���( -X�H�q����ݭ�(��,���h��Ai���V޲P�3a(,�N%��"׍�z�]{0ӕ5��&�\�]M_)˳���������&�e�Y���C���.�����M�z�y�PR�%�x����o��]�e�ⶽy�J}�;o͓����}SW��p����h�\�=dN����Ģm���b�-�?I߯N�uv�/�|��!0Y�t�3)��?zیzGu
��BRD�'A-O����4��#c�C�� [�����{�B����ɣ����jd	��h�2E�c	ޅ��&��e5��{����5��f��'A���9��_��UJ0��^X�VJ!m��s:4�9Yn<�.uP ��r x�Y�l��X�f@�&�+0�3|�V�>��n0/��g�;���-��ϭ_<�Ë{/1�ƣM��3`k�y�!�6�}������X�F/���Wcbe���*���h��n��1])���r�w �U��^B��-b��LqF6d򟗝t
s����6u��C�/*Ζ��R�ޟ�j�t<'���'�_�u?��I�Z�|�j�hد�b���I�ɨ���t��}#F<�O�ů��z�
&Sߘ�'��)�
���_S!���^׳�ܳ�,=l"L>�1,8�w-�|�w�;S��zqf�Ȁ���>�1�1����Ua���r��M���A�|xq�9#ř��3�8����`�y26�OɘY}�ĭ���������xk�|���E���*e��q�}M��Y	�ug�k�Yqep������_X́��E|G���E����|q����~��'&9D��
*O�M&��C$�M��4KI@f�2T��p/��+��M��!#���ʇ�� ��D��Ӳ��'xHi�|iaRK��ץ��J�6Ą��L�p 6~�ᐷ~!�wn�7�>�M�s���E-�q�ڪ7��l��(�>��@q��ƾ�X �a�E����:�î���έ9��^��ߠ�+U8���֬a�j+���)���U���6w�8d����;J�߮h�'�F�-R��/�n�lhQ�J"��V������j|��c�&�c�g��!?Tا�����M=�Z��F�דd�%�A�>8�|q��Pi��N>!�Wl�A3��&��a�fՙ� �$/�ih���4/,�� �:�H3�t|�Ӥ[l���qX@`�0�V, .��%�ba�!V�&q��ΖB��)��Nt��8�@����"��fW3� �C��:�H�F6��MN0+�4z�&\ ���Q��u�����Q��ˑ�*�i��xu�=Y-����ei�t�-	�wPYb�.RV�d�.�r/�ީ�,���AHxLAF��`3^~�%�E��ME� U�s�|���v��c;�O�zJ�q���|@p���L�y����՘��;MB�{�{ͤ5��f�]��r���F��DH�u�ˮ&����#R����f)�ǲ�j��O�$1�߈y�J�gÂ��H�;���������Vl�۲oѧ �����&sr�|�#l���E�:s��*{���7�1uēC�`ɳz����t@[ �U��=g��a�^�m��G|ċ��ھa�{��9y@�
9>�:睙l�,��]s ��ЩEa��의NhmkN&:�J���"٪���([�4�C�n���n��=bx�;����\��(�����`_G$���2��(6'��0�`�2a���L��_���"�^�$ƈ��é��Z8Y�_9�%��|
w�y�o �xx]�^�a�*]��������Tq3W����ԑ�0��zI��]���b`�]޵T�ᚽ����d��juÃ��˭}ѫ�j��� �m���VhY�;!�y�[����[z���EW�׽�[�e+Z�
��~�9GmM�����͕i-�����eBӚ7��YE#~:nv��T�z
͕˺�.mιVV�����ڵ���ź�7�����x�.��D��霾�0�oX;��g�ww������ U�*���YRx�Ux���n;����팴գ�3G���z�������~���0$L��Q��=SV�W>�=k����=��K	��<p�K����I�������B��ߔx�X:Y�}�h��v�7�l�&���uOԍ%bI�l�O��|.2�?�IW�XQG�B�u�oqf�u�w�����jc�;L`�8,���/�ď�����jV�u�8Xd:�a�r�����f����uf���[�W܋�>?�UR&��S�@`����]�N���5"��I��4֑��%.��}>	(��3�\�ϴ��Q?�i��
A��������)S�̈E���v|��������j4�'����sm�������q���-��y���尉��!q�o;�΍!M1�<� �5GaA/��Ȃ��c�Nt/�g[h��+�?�yq;u�����[uN�'Ǥ�D�D� G�Y�["�y$�{�I���TM����M,_	(OzRs$�8�k	�1(Nq3���EOҢ�Z-ÓR�����;��8�ջ�qr;@3M��ē��c� �Є��9Y.��1��b�����T\
�0�ȒuG{�UZXlxV64EB    fa00    2500{���-��ʔ��9����%��~ӿ�x��us�{�Q�ŀ�|��fH�s�i��<윉��Su�ҍfO�� `K��bx:�Kmt\�~F����$㌆ZR�A;�l��f��v�|���un�4��	f$C�KO��nX���?Qf����6��_��G����洞�P������B6�2'䵼oq4hNX�)�*��am�o+6���&��l���~2�E��4m<��h������6�{�ϒ�7ȏ��(/��6G;-�`k݆�ǡ,�ɛ�Le�"��#��v|�=,���L����hh�;T�Czѻ�-"�rnт�.�O�:�}��u�J�+p'�y���W�5���O�:,����=u����a�@Ai�X�L�׍��LC?y$@}Ys�����O�L-�0��p��w��;���o�RQ�P�k:46f�D�	������c�z��'��F�X\��r'SLL�<��;C�<��G��H�@F��y���̨=��l���;�,1?�\D2��Z��<��8<,nU�Y�\�7 �BrȲC�I���Fy�ml�x������
�Y�2�� �����g�yQ��Fx1$����O�`�H����%x����w��`>�����7k�zo���;�-ɕ�r0/Od�C�L�ڞf ��U�4�� ���j9.K������z���b������G�>o�m�h�𞜷X�zq2����S�0!�p�\{��D��S
�7��=�Oe�����8��^
ͧ�WD=9�߃���<IAT��h�"@�f��r����q�.�=���d�+0^V���$����������f�NL�����^d��t^�u����9�M4���h���L��"(+�#���@�"��У~��.�3��+�+_�+�)_,RtӖ��&��<��Qs������|C���G&J
 �
��`Y���}������kg�Q���j:s�+��rJ�����|Rrk�fxk�X��������%�e�F��L��}���	ь��"�?�ɫ6���>U��
�02��g�`��y�<QJ�������B��)<sk�![�q#*�'#�l]0l��x4=����)�t���Y]!��r���P���z��(.�� ��h����꼳!=�D��\�辻�`zQ�K)��P����M>	�h�1Ayi5�ճO�8lL^ ujVDPU ��X�7���y*���5e�m9�ҧ9>���u�/o=�� l$ׅ�R=���7تs3���xo�)o���YD�����=n�����Տ���>>q��ƩK�-� n��ڸP�����F�*=�[wm��՘`z@��c�$� ��:��q�DoX�Q;��nJS¿�mSz`���`��w@�T���SAF:N��Q��ne?�����W�+XIߩC����4��*A9��%t��=��0�	��D�[�'��-~�R�i��,-c�b����WƆ�ܑSշ�o��8X��?I��e���+�A㓩j�r�����9�:�7���m�G@��3�DV�U?R�����Wpc���s1�;�d7x+��(��S]�N���d���̗�l��y'�s�	�mb������m\�P�a�x�b�Z�Vι���莻�Y�����,u���(�B�u��JJe�n`����O?�W\���t�!�A$��<�3IX�@9�55gϚH^���R��m�x�x�+�R��yw0����(^�����0�~�$���z ��B�sF(�g���,j��p~���`����[��
b���7���ǰ����.�?.���3Vw>s�C��I�����YEcMT;w�NG�Z�5A�ī�5��o_��+��K㩏=�BFڗ��[����/G�Ӷ�4E������_]�S��'��#5���/�՘R�n#��|�!Qg�w5�i���p��%���b�F�;,�fkf�ک��g����רS�"�Vm�]�����"	�h�����	"�w<�Q�@�(����:��LP�w�M��D�����t/N�,7M��s�3�h�-1FʇОE�'�:�1#t��6�R��e���o��'��tGr	>�#� *����cn*��l):�U;�iU�{շ�l"�AO�� ػr@d�90#
�ߔ~��Quc�&���+rU���j`5�&��$��ql-[�}�P����EwǨO�ߩ��I�z�ƣo〞
T�85t�����3�>뾽
q*�ڊ=C��\��)��=�0o�R6��Ϫ�z}���^on�@��;m��
�^Y\�?�  ��ښ�S�t�BށĠ�?�8A��^To��U��s�j��8Pts�&1�*W�����;����ڌ���	ԣe�݁܄{� dg�(v�H�z-��?Q������d���K�@n��ᢲ�#ě=���r��x�)f_���.]�Gݢ���ڂ��i���%���pش �O��4B@\U*:6�A�1��YTǣ���5�[�Y�^vA�^k��z���k *7���
��2��m�p��1�
T*r)a����|q�DX�Ӫ$=�*�z`�L�ӣͷ���]�B�t=���.o#�w�܎�G�n��ԉ7�ҽ&�J���(�D�T$".�p��]�-���^��N�%d�w�Rv�$Jm��׾�aF�&�W���J�|Q&�=IuT�B�0jO�I����1O,�y
R���%��<�i��� P^#�K�����3�ìp�Z��G�3ܛ�X:o�A�B��?����]�Y� ���HV�Vu��
�|rӈ r����3�+�$c}�����Iu��H����e�༪q+^�vK妗�v�L�����c𯲈��ʓ]�.|�5'dC�9�sO�$����Z(����(�v���\����P2(65y2�y�%�s%�����Ȼ��q���6�C<
��.����w���Ÿ��!)�d�1-פ���I��/����mP��5ƱW��-K�<ec�/
��)����/�������|�jO![���$˴�ď7����
���U�	
fr[��E��4ӻ��":i�`�!ĎbV[}�;�)B�!�)�@����T����+�{���d$18@n:��64M�dt�L���%R�>�:�z	ak]E���L�"�}&���������ce2pdY��^P��4o������Q���p ƭ���K����j���BXD⨀��V�j�!|M���UW��C����RQo�}��p�mn]_X��b�t�?tHA+IE]3q�>;�;R�?xvŔ1��jB���������k���鮕F��
5�����h�sA+�?��۸_��	NK��N}��X�,1�8��o���R����~քŀV��\f�8�t���͍{���N.�ÏaK;=��-�9`Mqc�,�ߦ�D��`z��h��=��Wy�����ŒE@f�F|뽏���ky���ͱ��*a��h5�]����M����8��d�e������U����죮��b�A�ScL�Λ��j�+��=%�&�~��Ju�mH��B9�_����Z$��,Ԓ��ԎbV�v]t�p�frT�U��!�}�-�@�$\b�u���}��'ϼ�w2�>��mJ�#���q�n�@��;�@e��	�q-��	�@��-��-����QfP�e9E~��?�v⢺BĠ�'!,G�ֿ訷���Z�'ݑ|ۖ� �o^��b�»�h���SR[�g���i#Bi��#��(3�;9MǘL��R���ϣ�%(��ס#u@wo���6�=�Eq!���
��XG�V���O�:JxL�-�e�g�k&�A촐
h޷�c�>z=I��y�ҫF� nUxE��!�[\�N������3$��ςQe��gQ�x������U
��۩�\7E��Q(!����qE�_��Ѝ-�D��񳳩���&7��]{�)���Kq��gr,��5��I!H�|��%g��MR%,\mTB��ޡU��,c'E�]�z/��W��[Δx���c�y�J����=>oe�m��ZRLY�噥g�%��9,g�9�a'Y+�?!hν3��:��s����N�WBnkj�a��T�����������xײ���`�d�{V�M]�a���&6C�8�7����U
���t1���;t��`5�Z����W����vs�x�YߔW-!����1��Q�˕�L(U�r3	L}�H	đ��)֦�F�Ζ�k>���E��0晦.?��i; 1��[����U��avF��9!t�T�?�܄���g�l(���F����jw�ev2��h�\�L�J�7ɟ%��K��Lu��l��n��)�a�9���ʹY�)W̘��np��Mv���y*��܊:2���Do�;�W��GQ@!��vƦ���3'�^�Y��q˰ڃC�⸜@bUN��:$�2f�T^zO}�ݔ��&s�ݯ�R�T��7�y�K7�M�z�U�y(&_�ֵ|o�?.u��M�0Ajh�hεQ�1l]-eVT�i�f$R<b#-�P�����3�'�nW���6��	n��j��%&�He�/�h_Ԉs�6�q�'�z�7�˱p���80�^�^%Q��^I�����qL�MT�W=z����q��H�/�q_t��3�+μ��eF�8��ȝ���E�y��b����P���|4����VTF���b��rb�®�]�v����:B�w����-��%4_E�� �(1�{��專A��=��y�rhH�^MU����r[�5��^����FI6�������m숮��$�����Ų� �W��I�E�`x)�'�}�0�f�4�PY�[�;��%A�ګ���Ye ������?����^��BO��B�p6��}��p&F,�8Wy{S��ٛm^*W�q�����*a���Y�ƃ�վn�uUZ3�)����C3M�=����_�'�ZT.��vW��sc��(�Q�8� �:D�jY�32�.�s��Vus���M[~���x�S�\� !x�,�{���4cW�~<U��֓W��/xɲ��z�1��I���S��EfD'n�G/�a�����?4v�b���х��%B�;���ܾ��y��/{{����33�3�]���)�yV��$+��ICq{��VV�� D5�p�C�|XD�M��P#��ޛLۀ�
�W1!J��W2�s�r��;����zo�& qD]U<</M��w�g �R��F�Z�d F	<���W�������]n�:Zۅ��Ճ����6's��!z�U!� ��J"�|�v�s�����I�xg��[�������A�"����v*�_"�3�J�|a/cQꖱV.�(���2px���@����N�MU���H/;U:P�2�
�|%M(�S�Sr��f�HKA+�0�2�p�Kԡ1؍��ШDh�b�*L���7f�AKL�w"%c�%+��LEw���:|���m��xU1�M@�$.'\ܙ�b�����Wَ ���u�9^�Ed�^bؠ)R�'�L�z�ͽQk���8�W�ҫSZH�3� �P�߈Y�����ٳRq@! U���5��@ɽ֩���Ǫ[���gL�Ĭ�J�4�P	�I ���?Q4�@�D��nz���7&-�߮�G�>v�y)V.)�� ���ĥ�3�I�uB��W��Q�`SW��; ��*I;7���4�
�Q��@��=�R>s��P��G�a����bN��xC+\����M	r���KWx�m��@E�=���ʮ�k�C��:�<��H�
���i=�$�i��Ёg@��9��-��.xϸ�!%B��������
��[v3T������<��]E��*I
��3p�����:]�;K�j]�{ƵPf
��{j��2�
�rd�p��5!!�o�7f$
��y]�1�c�ןX�T���%j��w-��h]M�/�Bf|	�j����_�_�b��/�`�Q��ߌ.�����]� ��)�����)[W;��j���I��m��k90���%X����d�a���Wq���@!��Z	E�\;��J��ݥ0Wm�SlQ���=L皧��I��VU���ͨ�?&IZ��p��&<N9���hx�"N*�+����-j�����/��9�ᷴϡ��ʹ�$�z��af���׌�@��55cɔ]"?g�j|���,����;�w�)��xa��dE{�)�Y��tx� ��	�r_9x!Ft		��I��>&MI`#	����a� =�p��Z'��iT�����kr����s�TH��R�zb�pZ)vau����x�,㞌^�-k���_�󚰣����E�K������@����8�>ͳ���>k�ի�����$�"o狉��"�Gs����[���xkY��b���9ebc�d��Aq!N���4l���G*?k(��q��+�%ݾ�'x���
��!��s�
h��� 5ԯ�h�-�*��e�4��;M
/aե=�A{&a�*lz�51Q�c�tp:֨�g�'��?y�Z�%Z�m9���_�])��E&.��G���޺�Zm)#��>:t��Me��G��]�<si')eOXd��ڒ��t�}~�TWm����-J�8Ԡ��|�˖!�ŵa��@4Q�->�}4$��IJ��K�K=���g�J܇5pJ�z�ag�r�V"���^ő�sE8&��L��'�b�z�f��w:r/-%����3�N� �,��-x����b iİM8�5�_C���:p2��9U�2�=/����������B�zw�[��)���ը��n2av�c��K�u�IT{s�2�U��=5��s�7���E�A�	����_�r���	�zs�Oڗ:����jj��� ���Y)�����
]��%�[�#kY�&�r�[�T���NM�*����������~�"�:#���@Q�]�)�L6*���=�VT��+4��'��}�C<Z|�y}�I��J '����n� Z����������7�6ѯt;8"u��Kg�� u��J��B
o��YPG2g��>��Ó7V�mܟu�JF
�Ʒ�1V?jxq&}�q$ĿG�|�~���M��nH%�'�b?��y8�߿ˏ?�jU3�d94�>f��������5��n��Zg]z��K6w�o�Y�tG�,	��7���ݱ8�k�ep`<7�ޱ"�e3���<�&��4�魯
�w�2~��1�#�G��s�^?o��!l� ����U�\P��brH�h��o��G�J��I{�r���I'��^Ș��MXkQ�f��������"��w�-��ڊ�tO��B9��df��L��"�I'y������
>��,���g���T�1�+ۜ�I�6�Ey��l�5GC����@S�d��Qf�{,)׈��&^$(?T�sh�����h��oL���ޟ��>��
T��{�i'��q�5a�<}=�t���촊�a-8J����t���p5�I�Cg��k�Gi|e� �L�E��8���G����m�<��F�-��?>���`�1�^�"}���6B��su�����OH�7W�i��H3%z��B���4Q'8k�/� ������9���:�9��_��b�_7F�1M#�: =)�� ����������C[b����( Q�*�ȸ��-Pr��b?^��Z�+�0�
ܥ��A�$�\#&5hn��ḠS|!(Ra�>57R�aO^�4E��Ï`Sp ��kn���f}���.�2&�`�dV���b�Ӗ�t����y1���#o#�x[+�	_�Ȱ���s�y�URւ���ⲏv��W���O84;wW#��8 ���3^����(�g�h+��,�覯��j��Ó���H��i�]�@6SVW�JNә��^�����I����lǧ"S~T��tD|�SM�l͈��r������O͖� �����Ph1����H60] �&�M�,��S��|��/Da?�%��pp���p��cj�;�#�-��=A�h2v�-.����������҆/�T�%٣�w�A�J��'�&��}������t{W�:�uf�2}>��v��F�4X8���J��N|*�t��с���J���OR��@�[3?��R �����5�����`�Ъ�kv��B:���1 ^% ?5p�&w�����j����|�`e�|0x�t�׸K�D�������B�?��"�S
e_�^Jn��է�s��  ����Y.�X7���ޅ?��8)�q/L�-wh��%��?t��(>�)��I5DEL��	 M�M\kl_�z
۹�C���H��t>��S��y�7D�baċX@K�k6�F*�j��WUA�<&ٷ_�Y�����S�ٽ��g`��LI��Y��q�����}e��r�󨇱4P�G(����-��h�Wٟ���GsQ�`|+�K#��'F�S_Y�NM���>LAN<���y=�� �[���L�k�S�o��a�TMj���# ��p�
A��A��;���Uu�Օ��Z�x2�{��~7�*���!E̱4jUj�k�/�7crc�k4�i���e�W�"t0J���:��\8�K~|Ոc�!ffE���Iy�4���>mG���g�������eXtc%���x�3�;��o(d��y@�����7�*��{�ZD<�O�_!�I����@}(l��]�Tn�	N�V������y^���xP�~�k�ӝH��a�<� �³>G�po�$
w���y`�g66د���8�eu����"�'�69|.P|׳�I@_{ZM�)�MP����Q�s�%�D�������O�?��6����E� �3�� 4�f�DdD_�&6348
*YOݚ���VCTW��P��C�Yb���Lv��tZ�� ��}�h���=_b�Ə�1-�3���{�(s�WUzQSʻ�8�P\�|�hg����ޝ���T:�y'q���Œ�g,��� ��e�[$��8��؅z��|	���kh���u�ƚw@�Y�}-a��]A�>D�Q� ��D����i�W+}�ʠ�>		���*Z����F?��
��'"����E�,������K��e�/ۯބRJҠ�z��~�-޲��c�)�S�ف��H��T,wٺ�Z���$ؠC?t̌eU�z@���ܡ��+8\ �@_ �1Rk{$j"&[9]����]6c��c%u��4L�H���=70�h�N�|0���@�?��AȪ uSt�>�b~
�o�b���7\��0j}?$1I0^~1�6|�����@E��y1rQ�d+�Tp	*��t�ȁ�����`����X��D5��-5�.&�Oz�7I���y��sԟy�/�1������P���G���������HH���H�/�XlxV64EB    fa00    21e0�d����_ױ	�����O͐z�c,=�l^�A_�p}ǉ,G\A��i�ws1�N��L���wU����<Vy��
�)�{�3��S%��I�4�l�����̵��{��Z��-��#�sk"���5��}Q�����O�#ݗ��ಉn��@�԰blf��;�T ��"Y����u{P�x2ʵ�E�=�6�j[!�&_��s���W>���+R�h;�F�U�İ��?eۥa������h�Ф�{���Щ�v�E%���C�h�R����Oǣ�����k����VcA�З��럂���"@φs5;/+��@�[u�aJ��jEF�z�@�Ѕ���W�� �[�8Z���c�bihe.ܩ|�˭[̆q��,�J�e��H����ӊ�7�K�{�mn1Eg�����$K���Z���#]R�D)(��L ��nƿ8X��7�e����	���;���lu�;�ͱ;j��/��I$N:	=�������?k=9w�4�f�D������|�A����������{9fc緕��,ȓdH�����tىo6�!.eL�
ш�����6�:"�MA��${*�W�.P_�,�nh#5"��l����~5]MyH�Ѥ��O�	2���Ζv���f{p�a=l>���?���g'5�%qz��|T�������<�g�Ν�L���OWӲ�&T��2�6C�,O�tz��n�Lix4��	H[;��/��ľ��-4$�\fr���dΦ��[dPkAUQ?d�~�669�GNw�(p!;d�	N���>քuJ�����2щB��I�J���g�k��B���.,��oSw�����dcrA�H�u���.�~��Q���L]pQ�˵EhYm��~2�0��:n���U�͈5j	3k�,؟|M��tӗ3t�p�$7W5m��y�-z�"<�-wF:}�D[����e�a�v1���r�B�h�G����Z߫��P�D||�8z=l�C���ڍ�v�8ç>ɶ_m�A1#Q$U~�|g�%���vݙe�\��~�Lx��;9��Y�yW�^&�ٓ<-��_-�T.�B��Naa\Ø�tN��/9Y#�E��G����Aj�==�y�d$'��	�g^�/7��3cC��H��nM��f�B��-i��.���
PI��*���C0�9�8��%�#Sv޾��]RV3+�|&�it�=��<���,���� H੿k�(0~���@|����ZR+P�>Y��n!��֚�U�t�����z
1 �v	̂���0�58��;�cM�M�^ΟCÄ��M�{�.���H�1d���n���m�NQ:����2(#�XA�@��k����!b%�]7ލ�H_��UOe#Ј�9nH�Z��L�C�Xa��u ؤ�ג]`>A������U��-!���ʓ��ge$��RE#C���k�V��F��e�j��O�c��P��:Ĥ�iڹ������_�e0��&�:^T\QW�_���T�$���^���է��Wb�S��ȑN�ŋ���AX��wQHSm�q��ʥ'�{�z�9E|�Pg����X�ϲ��l�XQ�i�@6�z��'2�TTV�� "a0����F,�^�m8"hZ*��ygf%��O@��a�6`������=�x�1��g�b1�����oY!��t���-ҙ�rlطn�J��*��|vå�-�8k�9�6S'jA;�/��X�<?�[A��ǈ�ws`L0�6@F��7�@�]��>Y퟈��v̧��_��a^��ro{"� �'�L�K�����iE��<r,��w��<Y�`�/Ff߀����SMgw����a��C`wgpþ���2��#+�zA�n�u9��_�I�e^�K�/D;h���|����ȢA&G�d!a�d�/+&������9DV��u��2�-f���� `���d#��:(g�'��+�#騂�X��k����gyC@�
e�'S�Ugɩ���y%�k+p�
�H���ŉg_8j-��.4�+�3^�q�P�
:�ȷ�b�2�d'�O��P0%�Y�O�Mb�K=V��h�[J�/�|�ff�	8u����\����o���7��9�>�=��:"�;ڏE�.r�%�Z�F.},�MW�m�����#��>�2S��E�|�0`��L.	LAGx�,Ȕ��X|(��ˬ��iP�F�����AĒ�ڇg'��Ύs]�'������ա��}�Ak=Gg?�g�C�Roj�"��c*�M�g����An;�j������a�w���E|�R�d]�1���?���,�m�Pn@+`Ck������XGE�K	FJ����[P��,��^�Af�4T딷��*3��)�-�=L���0Tv�0�)���94�MJ�;��(l��(K�0�ވ
��bCD�B�/�Ң�w�˗�Y��
w�-Ű��Y�S�9��"𑃃/�e��Xd�9�iUO>k;;_�ށs���ț��iJ��\���_*�<u�p�y��ԋ�}�iZ~�ڬ�(,��&ĤX��_��g;Z{j����[�n� ��]���`�����K���%T���,�x�Va3�5=���W?э ���\Q�Vb�Fk�lfRA�缚h�\����f�|��ݚ�[�ԧ���̭/��é��?�kٚ�ۼ&�>}�s>m���W���m�Z<!���&9�1iz!��1ܳ��/�e��}x��E�1�^�(p������
��i�4s�E�W'��;�/���{�]j	��kZ���vWw>"W�������jP�3�q���]�F$5���g�bז��\k���NnE�3jc��Mz�4p'uJ��J�*�z���nyt��"Ј��8�wKYw\�%ܹ�i�-�e��N;̫?��α�D���s���ز����+a�u���J�q"%�|�b ����Qed������(e�@U���`n�Ͱ�f̫������ �w���F�S�O�X<-�I��.��7G�B�yfF"������Fǣ�����2���O�h��� �4���{�;�[:;���>�:�����#�dU�a���3���6�vF#Y��hy�������ͬ)��=��WX�Oi����hv��hB������a~�]&�*)N��.��}Q�[Iq�"�b؛j�'8e{��-�z8/T����΂��}D��޾_����`)����R[���4�Kya�OV����?#��g��?�#��h;�K��w9�u�S�D�7vVU���"����W�!�K��@|e��F����@#��8�P�A�|m�,�m�h����������戒��0�e�yjxh�;*�`��@H��o���Qj����?��]��܌=���l@����O��P;y�M�3��Ք�]3�r-�ّo��:h/���!ܚP{:�O��-�E�w��J, 8�ۭ:�ц�_+�

tA��#�wϘ0��=���ߨT0E%������5�Cjl1���b\��oz0�)��$����=c���ԣP��؞� ��~�hHxqH�����'�qm���i���r|)~�`tP��B��4�Q5��V�u71��d(ڙ������茁.s��U�g�?ѡ+����έ{gƦjK4�h�C�7�m��&.���<��ۜq{c���`��+�
E_���/���$���"�8< w�t'L�$=9��#t�i�sGc��5_���ۺ�"�Fߚ���ۏ�P�H�+��_De\��2��ی�8�ż�$l�H��5�ʒt���˕.Az%��bDB���`��z�>��f� �be=�=Z	�Í��_�_#����m����U�w�gܲX(/���J������e޻$"I��;LעZU܈4�&sj쬏$b�^����y�lF5�)�ȓ�G����غ �؀,ͺwݫ����J��������%Վ�����nZ���mA@B�h�P#Sɪ�@�w����6$'v#���-�V����
?f��J$7�� �^Հ�!n�1��/���@>�SކȬU"G�'[��Q�]o�%��z<1��y/��p�ƙæwZ�̓�p��"���Yw�D^�0�%�½:<�C'�������P,r
�wG�e��$~�ݱ�|�ԗ���`��}H$6	�x�B,��%ȗU����	�Ⅱ�ss	���ǁ�쩒xǩGǿ��&��lg0��5����L?��N@H��X8ݛH$���H���I���\��3ƿ?�{�}*�E�y������ˑ��Q������L�Q|S
�Z�7��e�v{�Oʐi��ޞ6 ��)e���.H1��R����4\�{�I�@X���"w�N�@������c��
�2�p����v��
<�Qv�DRz�������Μ���d��6X�;wd 6���Z��6���P(�~l-��i8w�"VX[�UQx5kȴ���"���N�\�s�s����-2I�̏=�C�Yw=T�*�&m�?�w!�ڬ��j���ъg��kw��h�F��A��
���l��GA@�~8�[f�U6K�<���t�����͋�ơ�3t1@����iQ��������L�o�G7\�Fs�I�}�=�GGgM�E�q���#�֖�J������J��Эgeb�ϲO\�)�=^>Z-���]��}�"�I�ZIh��E�8�f(9��lD��:IP'8��c�O<����8���ҙF����B�G�L��FMK ܑ|'?�ѩA�1�^Q��a��ׁ�?u}N[1����z)m�r�R6/ɨDie��BS�9 y���=���
F�F��Z��y�79X��OO��3���Q�[}����d#Ǿ(-~�u<���UóQ��H�X.Y��[[�0ة���3&21�{�gj#`,�Y}|��e��[j��l.Ca/
e����	^���H��݀%k3�� #�����/=rY�pC����4v��㧁����q"8�t3�6�=~8����ʀ�]m��e��pr>�{|��R`��� q�~�؟M�Gd܏��]�z����=Ed
�z<�����2n5�UE�a��P+�>���7E��}�yo�1��$�˫���y�З�0����1��l�W\��|�^����)�ƭ�9�M(_�iݴu� Qg��(��,?ݝ�*P֘b�۹#���@8�(�7���y����%�j�V��.��]��?8F�WM��xGᓤ��IǓ�[#~_�_ H�R�=\u<(�YJ��9|;�}uVa8�f�W3�wо�y-`SS
���X����D�(��Y��K��A[�uլB|�;�,�ia|}�@��o�R���~ؗ�mT��*6�5ԧ�q��l`���]�����.��M;�dB�%�����nU����2	v�e+��w�;��6��J��6@���+qV\����xB<	��o�J�!9��BO�J�7RPkN�����{jO�a�����2p���	)O��j`H�Xz�'<�+}�+8���J*�H�ݙ�v��^�oq�@��@]�q��9�I$5_{Gz}��Wm�C� �ݴ�%}:e��X�8ҼGy�V��w�N�$"�<w�&EduǍ�fo�kd�y�UXrpk��fC.�'��۴c5�������H���Έcvh�٧g�A<�5G�3�B�q��,��pG��%����Ⱥ j�qC��L�|��d
��kbNe���1��~[.{q#��q�F�\jsÖ,�#�-N϶['57e�0���
\iq���b���������y.4M㢳$�k�%��⿲bv�Tx�c^6(��^�W�k�`LXm��O��b�����w����Mզf{��3]e�=Ƹ�����U��� �38��/��i���3:�-���}U������Z�*x�nf����Ν�_��ϲ|�䧐i�j����nB��HB�t4U�1--`����caB^ju@!!ڱ˃�i��&��u�z��t���`��kFv�!�0Bךs�}��^{H��l)�g�Ԧ��W��H�`*7+�+��g,g3�t�R-6�, D�@����
%��i��{8#�h/K~��?�(�s%r;
{���~�?]>��6v��Q�ޜ�`�x-��
�hO��s��l�>8��B+��@ ��T2�:�Z��{'�&�ԇ�q���5g�ٌ�fV%,ܚm���
#�&�s���h�zn��`��b�3ǔn�ZA�@�:�|ހ�I`�}y�τ`��;Ё
W���.�Gn�L2H-z.��N�t_�}���rm�5
�Q����vn
U��V,A�������_�m6w��h�Sb%����6Ht�t�s[��D�������G���u�<J�^t��mͲb�g1(P���TR��t���;�#<8�9x@���`*���1;3W�O�����%v՚"7����һj��8 )���@���7Imp/��{Z}O�#ڋ6��M���Vs�yt5��r&��zv&1ꀰH���a԰�*�F�,�����^����I��8��BkDmU�--�7�mr�QD`���,t!��s�4��M��ty�B�c2-������9��O�}���頲�A�w)7����U��۴���N��7��Fض䜈�-^���� ��y�QΧt?�>�,�KM�
c�]��[_a�~04�Uu��r�	2�~�4S�x��d+`Hgv2���Hq�Pd⛌�eby��ipf5
͌f�s&��s;{M_�rߕ��E+�������g��~D���M>0��@�R��r4ʳ�A���o�_G���dŰ{N&@Y���G����vB�_�����b}�2���6'-ټ
;(��{�%t�V	L݀���U�p:`e����[R��M�Q�����l���h{����R2�S�NK���6��&���d��s����UG�E%�^�"��fTk���|��� ��ۼG�P��X�'�Dǽ�3~#L�T���ɩw"�E�c�_�T;�8<^�őM�F o.���ʕE`�u�h����SD�fvܑ6J�	����1��ӝ�����g��U����ƀ!ybFP�`7�U`Yڴ'U[)؜���{�l;��D#n>��x�W�:R���E9*�L{��j.�a��󎧝�U~��Y��m�e�<*��-�~&����l��x�����/Z�ؚ1[X1�'>H����Գ#S��dF��� ��/�lߒl�"�qU|�I�B�f�����,Sځ�:D;߁+�脃���)���<.@3��'	�6��t`�M���@��IF��r�>pÔ��#{IT��7���3�8E7t}�ԪPW���b�7�ɲ�q�����z+%BqZ ���ݡ�eW%N�:��3�>�ҽ��hLiTQ�oR�����g�6х��R6G�
�*1��ף�M��Vaܥ�����K囻?�6ճ�S�
��!~P���p��i��LO�->'fi3n��R'�"=�[.'5��Ϋ#"�buP�nA��v�e6�j�xY�>NYs"��_��v�v���(�v֕�w �ķ�C7wiS��K2��Xz1�!�S'$�PZ�`_]P/��]q���y��F|�E��3IP��L��-i��X�t��z���|:Ĕ~n�]Ц�� t��U��L�E�O[gC-��t:�k<��S[��&�W3��,����.�6��)%��X��Q��_��<8*��Z���벖��`��wB��7��~`3�w,��FL�lV�3>z�@�6�I�N(�[ .�8|{5X��A�M�x1��X
WǍ��O��j�7�z�p.�.BK}#��J�o��/��hH�pce�_�skl{�[�B3~Ė�{H݋�R^q��|���z���)p�B۳�ID��ނ�f�Rֳ�)*��8>�h��:e�����8�/(������)���D<Zj�%�+h��&�~�9Rf[��3��Y��%�EN&�LNƆ-�t�ե�$��aN����IF���ƣ5��<�?V6n��Ӣ�1:�J�+��3d{v�:0w�����ʪz�\<�m}3@�X��U�jH�l��g4�"�]Lg�wP�ܶ�x�u	��\�� W�.h����+��6e<�LeS�E,�!�<jEA�S��}BsТ0j�_�� a�$RY�A����4%F-tA�2Db�}��/�2:�O[h7���Ee�uK{����dq�s���.cͧp���Fԧ��.*� ̂�rY� d�����b�3���.�r���h��}�m�%��[��8�,����3G��=PG@Xk��jh;#��r�vc�AQ&<�]1c_�O�}M�y���t>��D/����i���B�:~C�ӭ�ǡw�p�
�"r͠�
&���ل�G:�����L�Zp��Ss���=��z����v"�^A�)�
��)��@s��l�9[< &U���]�W�L]㱙��s]���Q8GF�9�TTH�g�;h*���\��c��BI0�g�}:i�Q"o���-��֔�E�_?f�f�NB������Cer��Ő�0���M�o����6�c!��)��C�-3w��/��2��CµWaF��?�%vU��ˍ2����*���k�<�t4�=��C=�N*��Ȟ�P�p�B��D/!�k�$��Nm�X�B���Wf�f���4����6W���x�HXlxV64EB    fa00    2560��s��(x�a�k{��H�!�A_�v�����������vj��8�x�J�UTfV��b[��2� �T�T
�����a4D9a�F���$�mq�巋-r˸��̟�s�/���L��]��2= t��^�A�]�%o�'I���	Xd8�'{�5[|R`�b�[��5H������nV�~�̼ˢ��15�m2hp ]�y
��&f�Ec�,=�VAx��*��y_^K�0�W|�N�o9?�'-oV�£�ӫ�4������K8�YM?(޹�O:�*3	� 9m��x�I�&��<e��3�k����֭dOL���~�t6l��.��2�m�ք��3�MR�~��΋�&�݁g�`uQp�*x{N�>�tc,����z����f'�4ð'�c�)&{��ת2Y}��'N�n.�${�Ȱ���aFp8�U�^a��}�����n�I@T�$\d��B���SZB���cU!�����]�vuW�qWڈ<��\���)/��L�oe�ȳ��;�m��p����L�z��8J�eN��R44<�kW�y�a"U����w�H�JQz��%��n:����V��Jll���hk��۵=��(%X���qx�<�wB�&��h-�
]��K8ػW�]���D?������{�Ӧ{#ِ���U�y,�9��'#�w�&룄��F�O�m���&c�HY���sOM��w�h91s�h��c/:O�x�le�%��:�Bf�0��"z�R��:�%�Q�h� 4�0��0���������	��Jd��ThX�N�z��ىNH5a��a2k�J��Re� {6��0B�tNlo�3�9��V����q���>�G�K��-�'17�ɑu����%v�x?��m����y ��W�p���vH�[�Mu����[P�M��
?�<pqU�PV��Љ��S�э5J��:�z��l#�-�@a%K���ϟ�+�xp�\u)N��,Bo��Hڄ�>����w�#��;;�����`_<yZd��֙��N*���B�|c[�p���~�]n��k��EH9����&����L#���`��&���M0<Ρ��E5�a`.۬K����)z֠����b|��z	��A��Q��V�~����|M#��e�����oo�b�t�ŷ�,w��nP���E��5燭��9�&�g&��DnҚ3��=�~D��V���%��Ǵ���+���� 	����Z�����W��ږ@m�֤�XN7kK��h��P�:৛����Ƀ)�)6.v-�]�8H���J#�а�0�խ~���9"��*@��e�z ��m���֑���X7��y~@��2z�7W�T��G���S|�5��
�_%b��g
u�z�����4tM�R�c����m�
ox��u�iKH�橋��m5-�I!��z�2���� O$4�#�
���HP"�q�m���y�Nqa�����-�amJqZt,zjR��JB9'�>9uܫkVT���|f&�|nP0s��h���_��=�����_�ϯ�9����cM��d�����۠�w�x��F��QćMk�
�ow����FPk�]���
����W|��:%z�i�ᓎxe����{��ђS�ڏ��N����x��v��aqN���h�%��є3�$�5��h�b���f�g�	�(8�W�^1 s�ǬJ��e�+{�-b�\��9����\�#�l�n�iN)�C��� 	G�Ɂh\����y�:�|"��޼�}�Y�B��[��\@d��]
䬹>7 �>�*��~k�2KK�>���.�r��e��4f0_�L��3/����'X��nOѩ�w
���CU��M�|sc$��=â���>jʟ�S.W�}�ޏV@�p1a֙y-���^@��S�������}%���OM���~�͕��#�l:����}�T�뺒Ir�C�}�a{������Ȫ�c�j�	ؓ�
��N���0�O�򋭻����瘬��5L�k��=uk��G�7���n��5�J���tV �%8p�y�`���et�[� �B��A�2�k�W�r�㑽*S�����\�y�a�Z�SM�0��R� ��	�h ?p��'Vb5 m�M¾���0��lވ�!�x5����vuC�c�������I��27��;���Ƥ����"�5�5[7Ea�m�F�(����է�5�ſ�9�	�;��^ ��'�&�P)���&`��+��D�9���1J&�x/�E�"z�;^���0"�+��C�p*\�U�v��c��έFZ���W��g\��M��>P����[4�WU�d���ǆ
�M����S)���ī��	�ȳ�2�RA�Z�M��;�toP�j�P�<�N͞�s�p嵁
��1/��{ZA��'Mk0U��7*�4^R�o]3�ݺn��m���z�5ҫ�����M#G��J#�����@��v�~��L�A�p�N��.9&б� 3����2���hJ��C�>%{Bx��l��v$�I�8�5�����Jdd���W-��*�Ãv��^vC����QrG����xp`���6����"���ݼ�:�۟�c�JZ}IR�|�'�b5b�B�BF�xJG���	�����I*��cϴW�֔��T{`%�R����-�����;��c���$of����س��dY	�R�%�g���4��D4X�C镦�j��"2o2�u��'Ş҃X]�LHk��VA#�*�D?�]ϰ}*�-?8l�2�GޒIZ�x���������p�L��_1(�����}���䯝�(�t��wcbr�����!�S�v�<��q�^�q���T�Y2�9�Dd���>�^S�c!��R����!�K��vϦ�n��,�8񳿼��e��R�����������<�y�X濧�D�xh�lAJ�]�
ڱ!�n��~��v��$Q�]{�>�p��w{ܭ��%���*���/�N��s�F�z`��N���()�X���#c7
��^��p:�%�lu�z�4V�z�E��#*j� ��C%�T$�Mܺ/[;�CcL����Z`��	��'��څ?u�|�T4����{_3�L&�{D�B����%�$���㌈H8�U��42����+�^�X��!cM��f�l2�B:c�r�Gu �?��E2m�vn���1Ŝ�Wr����9��Ε#r��W�s�$Y��6CC�rF# �2�#T�����y��F��f�e��[�f� �I�{�x;j'�"�㴫V�hBs:cؔ�z	����bL��8?���65q��n �? k�₽�X��|�/�jt��!��gq�w�B��ݸ&���`j�=�︼|$J˩�5��黩���ʴZg,Äp�I��wm�ND�}�c�%���nГO�-]�
9ֽ-�Yx~��o�G��H����AR�O�2f�7�
?�����(��9�f���H��auF�(ѥ_Mp�ݍ|f��0�y��ӫ_�ٓǝ�%jH��oN�<z�m������(`Ï�K@U
��[f�7��i>�����z��V��G<�+JV7c��>��Y���}��
���"��*+r�X�"1��2�Z:���@�OJ���ߓ��h�9�=D��Bx��S_b�'~�^��g׿k�3�*�!m�H��h���X|Q'��20a�~N�,LȐ�rCM��:S�9�"����@�d�*�+����*�ԓ㏟�5m���31�=�>;�1����.�	�ȧ4!�"���9��V�S���3�<i4]"��fW����m��8��v��N�߈L�@K�݅?h_����Q��ދ�i�!	�k9 u��_'d�ǧ�%�@���Ã�[��މ �*��!��t�[	=�.Z�5@-��/dv�P�M;6�롿b(���@\[\����n$�N��!(�GQŚ��U��Ⱑ�o0�����PDw�ܠ�IŞ��u��'c�K�2K��ģ�B�����rn{)9��Sğެi���5%��~�2]��h�h��Rcs��,,��G��k�H�2�ʀ;�\I9g��	^�%��ž�oqx<�k�>�Ӯ&������lp,�FSn�IY���Ԗ٧��˄F��~����e���l,�-k�FL����v��gy�c���`{�'%��wWq9��)f�UX6c���`6F
�Nd�Г��V掅��,!����sX&���Y?"R�笓2��Y\���MZǵz�����t�ˑ��+�|[,���a�J��I�P��%9�D�ޝE�inϒ`ڌ#�7%�K�V�"��� $Y�h��DV�@\͢�.Z�&�z��X`��Ezź�br�X�q�>�܏�N������-NK��x���.}E��||o��z�[���ߖ�C� > ��,Rg��J����oN����'��f��4� $�(e�N��v<5�:yu�I��%p�(�RJ���u`Y���$�6��`�;fYI���vB+��8|W��ˍ��~�������7VP��4q(c_�c�k��O�����Ǆ%'Oa�u�֏�^ǿZ�/�=�N�	P ���,�<���q1��C��5�w�0ѓ��H���/3~46r�Wne���k$�1�"u���]�>������Ț�`9���@���p�oq�ȗ��u�"[*�%��(��^V}�X����b��~�M���m��r�;�1y�)m-�}�1�Й5�VT�cCV9&��f�{�=Zlq|p�o�K�:lGo���v̙Ks��Ce���_��&���ĵ�k�Ͱ/����I)|��B�Ϭ�5���H.2�7�h�IQ�"H0�VBd�X�����b{�wv����SMj��o�Q��p�]�0�G������ꉯ4ǫ������=r�|Cʪ�N��Z�>+t\�$*T!Z����2�����=L��s�PF�A����iƨ�ۈ�dy8��.`>������ٽ;�)��x"ɷS����y6�,�'�@����hp,͠#C`�9��w9T�ʛR����㌁���1
����Ç�\��KX�� ־�д���"m��>>ܗ�o<fc�T�p�x]c��\�^L-h�n�����ۀ"�&��t&�|?��:� �GdO����O|}̕��Z�+�#܀�|<�LN���b	���>0���Tu����N{��0c�1�ӳ!''ɬD��j��Y���X���x��i�� ��6 ���FR��Ⴙdk�Ǵ���gXE����)&�֦�����srSb�7�'F�wM�6zg�bW�/�/Z���w��7���{���f�Zh﹀#'A�Iqr�<A�;������Q���
g}�}#�kJ�t�P��z(�
���X7�'��s�cP���-�B��fE�cC�L;�PHg�1`gCk�A�i,΀��*ND�� �]����9$��r�g�_j�]�i�e�W#�$����%����.�?;������M�|���~�\+�t��q��j�����m�3�pJɾZA�i~�p��r
Su8���y��^ݬV�M�@M����o�?Y.�;쮓EPP�1�y�BV;��S��|*�r���qݽ��8K��U�4.��9�v�����Jo�]_d��y$B�4�fz��N��L�ځ�e�с���u��7v�vȊZ�?���u����/�w� ��I�G�a-ţlW�A���$�vRB ��q������)��e*�y�d�#��?���H�u��3-۸Q��9�b��~N�N��[/H\�1�X�$Kv �H�J�ly�>�*�54��Tq>��������[�jg\��r�,ή��AQg��dS�-G�2��O��+����/��YBG�����5� 3��s?��ɡqK9g�D�M-�����f�WS�Ӎ !'��aRg��yg�f�F��&xD��;��AC��u2ecL��|w�Mx�՜8X�s�]v�ݚ�Q8j["P�F�£���RG�Tw�����6�H�y���	��Ӫ1�_��[�����0��Y}2�,���v̎��7�3���V���B��R/Aِ�RWH�P�0�����I( `0s��[3��;J��݃��S�ƍL U�mB�m�X��h�t�n��f
6���X����J4C��w��}������t���t_?�R=�P��k:��IS�ա'!��K}�%XW����#���y�b�%����[r:������<i�Č�n���|N�u�W�f�����^�v�@�w9;j2+�&�mc�g`�<�̚���Y�Qp\�C��hd�Պ��=KP}���Gu0����XŎST䔆rVj�̩~�b�1=��`�_��l�~��.���������Y�5c���0�ͼt��Z�R#m�op����#OuR���_�.��-<�(�f��__v�����&����2tHj����;���z�ݱ�B��/*����w��/�&۟م��]Z5���X�٭����$)��ϗ��>6�s���`�O���%� �Z�}�ҏ���1����	���qĿݸ���XH��w�O5��9�<��,� з�� ��(�o�}~�>,K����№.gǑЎ<e���#�2i���#��C+ds�t-�b�~�2�G���1����zwq�2_�CeM�ޖz��|Ѿ�P�ۋ7��t��n���ܖ����cP�5���j����o�6slx
dKH�#��2g��_@jm���wk���E�:��� OUP��`�3Z��0w,d�.
�(��L�+)�q=�ӡu]��9(��eܘ��}1��Ul?�"0�xS��ᦋ�G�$��>�)�ĕ{fI5��-����d{Yk��rhFW�H�Kb������Zf���[�{���l	�*{��suͦ4(j��iY�\o�	3%`���N��})#�G��<fuI���]�ؿ�GڭxO1 H0M ��j�*��9J~V���!���`�|�dߛ����v�<4-�[;��q'�[�Y������t5w���=QAq8<�ގ�?`LH�h��>$�Ɨ��r\`�m������
Td��2���hyQ(ʣ3c�sZ�Oi�>��@EU�?I2�v!w>4�;~�1W�u�oY��Ld�k���qi	�ƿ�	
�0��=kk�$��e��4<���C��%���cl��/k6�H-V#{s�
��y�ᠪ��^��!�㵾��)��0o�b�����wʖG�^��-��xa�����"�x6)��x �����7|���X��޼�1��?����Y�n�Hˈru��z���iM�^�v��o?����L���.	�FCM=���ZD�K�T�<4?8,�@/\懦�?v����ƿ��A3�f�(lU1^l�>����Y��� ,Ez��R��1����>	�6V�̜�n0#l�z,�ovi������I��z%��K�-{Y*�f�$1y?*1���w�#y"�U
f�`1c_�,�Z�"[���g�R�ϒ�!��O������E��c/�m-�"Ƀ���� ��������:�������S�&Rj+��jd�[��jF���ګ=}q~%)��|�`��_���[�|M֧��b8L��
��pop��C��:�î���;�d�U�0b`�މe����1�$�~����׭Q�.��B��5�I;Ĺ�`�E7�������Uj��҉�
Gb��4�Ԍ�N�T����35CyS'���Eh�,�ߥH�]�dG�����s�8��Tڈ���!���Ȯwn��ux�hǹ��z�(c<�=v����W\���L|7V���?����x���h+	���� �zr��%�w0�_��9B��J&�K��,�:qZL���a((>�<��
����F�����v214Z_�J$���_�P�!���oT��9K�9c��C��漏V�)�R�w��9��7��
`,�R8�BR�����V�Y��gW�b嚵� =�?0�1O���vI�V�ŠGDə������v@t�����&����'yĂ�9\�!eD���y8��#k���5�Ȩ�����Z�aM+�Nfs�:�W�lȢ{hU��}ǲW/X$@�K|lm����W�G��N�NZ<���]5���]Q��ű�0gږޠ'��/��3GTe'��#�w䋜W�&
��K��&jv��9������>�D�~�SV��r>3��� gd����S�^�S�T$�?�YG'�LC�Wإй"-��t��l��X瑒�2Z)�@��d�s�}N�s{>����3��w�$lٹ�����ģ���g#[ ^X\�q�>��NJ�tR�'1�;q\��@t�oҴ*k<x#N�?���|mi���3KB�c$j�K�C������1`u[�C�"�%C�eD��x)d��<	H�Է�ua�|Yv�������t:��{���;/��Pk�����g��;���UI�P����x\��i�_�50�B���޿_��6���6놥uV>�:�Oϟo4�j9�{���`��@#��,G��6��_��Vr��᪈�/=�}T���\��̋O���X���	��|�!5D9�7�|)q��._�2�2Z���z?��k�LI�p�$��*�@L+l���UH"�K����b���7���Cק�6�������\jr�5��H�~eN3N��/I[_�-��Sʆ{�j�pלM�ls�;#�LҾ��-�h����T<���~�E��e4�����
m�ޙH����2��[��Sj<��If��@�<7�w q�1R�I�;
�N�T@ �h�ό�~��[���TC�oL��� 7�g)-+�D1�"��WQ6�$ӱ�:h�6rB���q�W߽d h{��g��7�F�T�Y/H���.@�Zͮ�Z�s�n�ɿ΂�臬g�+yIM��a��.�͢_�B-1�x��d׮���%��A%�*��)�w�%2�<�j��G��#�VsT�@�ty���<�W���Gn�+�
U��#V-T��'�b�߃�=ufK�垙���4�|M�z�6����Vk>�c�W�����Ҧ���ɴ]E�DC��#�k .��H�Id�J��2�mwY�:��1��G.�`�E�W�j��3E��~���7�̃�ms���z�j��b���}�1p���Xfu�e}Ϯ���m�r����^�nՔ#�F��_̶�M1�uq(�C����wgy X��g���y��8�|�tH��E������`L�|�j�S
L��п����M����T� ���
\���*%Y���y3�x>#dI$W�|`�C��j�\�`���-�5�aL� �� pw����[���d��G��ڀ0Lg�(���_��W�n�S�vL��]�0�S�>-�M���ݜ�$�V�
6�{�+������%E��CSR���Д��#-P��9���ɹ2� �6'v��ar����yco���I��������u�����#�#�,�.改�I')������5�*y�e����Ͱpi�6���XlxV64EB    fa00    2370�(3����«�M����7K Ĳ"�:p��@�lBFSM�k��P=�0�_H�$AM�.�g�<(�L�B�gET�*�6��h8�>/��*���N0J �`YG}���7$��'5�6����_��N�$1LB���e4�V�'����ǢԥFq��la���$#�֌zD���_N#� B�5���
!N�u5mr[�K7���uGi*u�Q*�*YѢ�j���1%��k]������៰�^Ue��Ij7���E�~��G�3D+���a�"���v&��^�)�/|�r����U�|��FR�(���=�V�\چ@�����ҟH�o,�+�	��Jm���*�3�h�T�i'L�H��x�:�2W�0Q �-#�O�!4�o8o����Yͨ�oz5
�[0�ˎ��[�w�)ݩ�ժ���o����(��ә��d�
A�G;�y�����*@m�R��o�|w�tJb��x5��6A�Vb|�؋2bǏr�c�����:#ةv�x�'(�:?�y	�#08�KQj��ь���0/��3���$
<�:]}�3�Ù~��n]j�<�|�~������Yër�~���h��Y�ť�cu�hqӸF��n��_��%��_�Z�,�p1w��1���e��l����=���N���~��ې�}�rp�p��x�����SM��I���s�8��vK��p)�B	���Md2S�u�e'�O�d2�siI� ʘ �3!���V�h����n��@�w3�|�g���1E�*���b�����p�"���B�){iǰR�'!A�s*8vnNyA�Z��d��y�OU�g�;�o�:3%�G3��Ĳ�D�Z�J]����c�ɡ��b^���y]y?~��:8�c�6�U��4+u0�V*۲�%���]8���xJ�ōg���q��ܑi����f��tܨ'���i���ዣ��w��vz�ڴ�s7�n���+H&8�}
�C���Џ�����LP�ud`�f�Ժ�ۮ��Z�
/��k��if$���� +x,���V�u~Q!�Մ��-�8�m�	��BKխ�<"ϴC�<6�@���,G�qE8x.?���qr�ӓ����3��]�1>����%5��C����=!s��RMU��?*�n�T���Kc���1HS�jL�[��1�a��;C��n��ѝ��P��l�ܞ��^�8.��wi|�(�9v8d��u>ʾ��Ц �Ԝ��E4� /ۉ�
�0t3Ȣh�B]ű����UɡʞM�_��*�Ï���V�ٮ(�T}��⣒NH���S1�;r� �m�{�(�^��B���K�Y�c�%�c��(�(�S���W
���Sn�H�ԹX�����o3�إ��dƄN��ia �$�^��N���Z��i��P��a��6gu���O���&<4��O5�;n ���g���[�pGLit4��6U�oQ�L���+&�>��&�H�z�����D4p���[\�вY�4��(6{�H2<;��KR4qB=�I�KR���0�D�W��yM&�s��(���ү;5Z� ��H&c;���P(��
���R��v��,���s:�a�L<v�G�/>��2~g���)�U���k�<ʘ�.��b6h�z�+f�%Ⰻ�Y��<Q\����ſ�ؾ�ؔ�5G@���9kyD`���1`
����d/V�+k0����<C�ט��ۈ3�g�fz�̸(�|G)C��U�!�&=����DJx�Z�l�,ӆ�Ĭ�@3.X���`��U|^�fd�~X�m_���M�%&i&�5�/W�8'�js\�a|��z�q���V|��I0��������R�1���Ro�V��.C�v.P*�D�t����7�L5��M �)�.�\�ƛ�?�$�"�\�OE�3�8Č�ML�#)#Ԝ[c Q��\�RhXF��o�e����a�������R����$%d�s�w��X ����KuC�EKLʸ�E8��E�6&����O �s4\F~��0*�:j�\�_��V��� ��n�A�7��,*�س WwN�B@�M�W�7�3s�
�*���dR���eXb��d��)}t�wЋ��Tq�rIK�GV�"�4t�º�Ǎ��T�B5|B�Yo9'�Y�r�(	+�?`z�.X��� t��[������$p��(�����mD�t6�蝈yG@��O��li��<|�s��|1�h�gsd�HqG��%[?Y�d�\�+����+��[�	gcG��'��c�"uW�a��?�:V��EگL`���Qf1?e��=]�9g������iYЌ�:��ݚ��gA�JmrJzE���Do�@׆�`���c���J�
3��GK��b�$n#w;���[
���C�?	@͜2��뜕Zҽ��3�^��d����_!�ϓ&�D=��MA���PL��?cF.�*���(!:%���?&������i�!�t��k��s�wj�XѤ>M�Q� �AI糴^YUcR�/NbGC�3d�8/��+��`Y�<�dY���$[�:�4U��S���toV����L��mE��1�Ž� ��N�I��Ϙ�w�k�4C��ݵd/S`�k�{x���P��M,���b����AZaS0h�-�e�|��b����5�4b@�T%Q ��3q��"�[���Z�C�1�u 1�-/m�&�@Sk1f	/���o^W�w�&�m k@ns�.�H^+7���ez��x�)���n����1���㨩]� u*�زB`���pA4�0����h~O2a0�b;����I4�q�n�~���,�D��۵l�d�2��-|T���]�Q�@;քY��Jt���F�LA��5e�m�{܂]���k��`�2N�?S��b�T`D������:�&c#��ٞ�]�4�GХ�@���X*���QqeJ9�8M�G�^�E}tl@+u&��S�:���})�����z+�*���;X����[b�r)W�s�b��*s�:����'�Mc��TnaK�)k̫L/L�iŪ���u���w�yWA�D]WU����R���P/:�Nc�=�Ep@�T?:[�p���������q��Ԃ)�t�&&�9 ���^=���6�n�����֎��B��w��'$Ig�����d0��D\")�,���v�E!q�*^	�Л[mN�=�DY=s��"�����Eҽȳ�5�f�o�ImV��c;�z���h�׮L�f�mf�x@F笜�Ճ�QI�[M!#��n����Dkj�^���o����##�A�X����@�ܒA�o�P�x�
��Ia����ԓv�j��{�d�ئ��6�$���;��Έ3ź�ȴ��!��w�ג4^*V���d�պ�e�}��}ic�3^0�����84��N&۪t_	u��p
�c�����\5��C?���W���PkeB���w�w��hK���Gz�}��+۶.�W�yzgD���&�\�LpZ\��N9=�9N.$�gm�w&L����Z�A.�}'r_sa+~��H��Ξn�!��mБ��㱅	�bf�]W9����5s���U#������|�Nc�>Aa�**�D�?�����~�IJ�ހ�^��ޡ����⛍aS��n���z��SIz*�ps��⸙��ZC��"�Cүa�����[��x<|4��9&���!p�34dƒ�W�EN�n�������
yXP��M�Y-��6��ah�L�	�z����St) ����ԧC�Cu�=��k|~g�H��S��g����kÊG_���	��{*A�Hў��>��t��\������,�<�WX������N��l4~:Ѧ���<�,�i+��{Ln�c�|tL�I�\|�;�Do��6��bc8��:N����jz��^s�AK��IH��#EU@���Yu)���s��˒���}?$`���eh:�$'���2ݾ�����߷�."�yn�gr5@�#���J�e���l�
5*O�B�>���)�'���jY�.d���q��ހ�	���6FP8û�@8�Q��@���LF��jz���S"�I��@�=�D�ޔ_+x,W���+4Y�|PE�9Pay�K�+7�4��Y��3�����dk��Ȫ�.��;��f]kl�t��	�nʲ�q�������UM��ns��-`�&�C�Ǉ�<��=X&�����Ɍ�Z����8_���̖���Sw�lmÙ� \�/-뽤� %�ej]=thq~e e��,�t���IP)�׬�Ղ��K��B�16=���̇�ڳ���'X��햆tz�J�;�����+�l�`�x1U�$q٠[ܳ��c�V�_K��s+� �m�T��\���Ǧ���]Ӊ��֎�k�k���_Q;��O���۸,2��=/�$��� ��G1�˗u|�h�f>�b��Ho�o����"\���Z���,¨�����קŧ>]g4�ÿ�˪��1��ٚiHq��-�æ���x�����Q�$J.GDT�K�;Hƃ
���K���\&�ӏI`�7V��xY�Sִ`��~�� 4�X[�E)��fa����^PY=@{3�pz��qӡؿ�� �)����z�5hmzfB��]�aH3�� b?�,���{s����<B�9����]!?t�4~U�M��TD�f�U�SQWSt�����r�n�K�S\/�y��{-ςr7O�ޮ��|*�n'AB}��ѳ$��0e{�8�qf�<1�� Ϲ�v�h�fN��9u����QÉ�6�����k�o�A�5�
�8;Ң!��������̫�*�.N�=�K�3�l������_�df���$>��3eO�NN��W�{\�E2*��#�%"��^n�e,O�02�;IL��F?���5C!y�Y��
>���~�1�M���_��B�EM�r:�?��x)���i�<u;�.H�"��(�1;������X/h��Q��������-���{ ��r6E!���yFX��\r=�$����i�YQ�ӣ��Y��u�`�W��v��7iOܖ�����Դ��Sc��AW4�cFg5¥��N���4
e^k� 3ɬ�Be�NԒy|߲���S��h��I��w-0h��aL�=�p�������	s�(
��_�.��hQ����>�#�2NI*;Y����2#���\EW zC�@����s�͇"��fy��=�X}P���	\�\��$7�"BV�����#�N�)���D��R�,,��|�P��Ka6Q6�g="�x
��g��q ���uND'���?5]�Mٔ���7�S^ %N��'m�1fT�#:�g~f��IH���זj�~N\�j5�d�wzb������6 ���4�2'*��o6��fl�\1e�,�Ӝ}8.����5#��§�3O�F�������d�y����Z�[aDf5.��nV�N1��Yy����� 6��:��EP??V1�B���+���S���# ܋6@�����G ���������G2��H�~ _��A����F�qVz5��Gj������Ɣ��	R5d�s��6���A���>h��x&s��.���&��I!�l�WA(hX�M]��w���70�uj&���/�廤��?x�J�)����n@����w5��j��'�u��'"J�y����~Q�M���U�K����-6o�ا6i�d����‶!��SO;H�/��H���ȅ�]�:�Ý�
F�4�O7��}w0��X-�#ma�ٌ���XT2A!�BkA���P��飄#ƻ�b�#�\-��VV�M������W��c֊y��wY=�m��7
���OA܄b*�}L�Ol��u�w�ϩ�*�]Gz�
t�z���ۋJ�La�o3i��F��Wv����;7��'���ea���џ@u�vӮ�=�>�<�z���d��J�C4ǖwqY��BL9�L �rT	n����Jg� ��ӣG5�Wk�.��s��ީ��y����ށ���}��^��Y1t�f��Bpc�_�������+(�r����w�l#��E��xW��V��m�*�;
ݯC��6���Y��E����M�/�n%-��:��@u��_pdu�_��x��)*s2�sˮ?�7���j�!%x�5�n]�
��o�uP�B�٪�M'�9
�q��l�ݦ����Hw�D�pjd����q�_L�����0m���t�Q���[�]Z}�T�'*�t9{�l��Rό NR_z�;��H(Z���M	�_�&Q_�9:bS�BD><p������N�O��MX��4�������^#��@�Qw�U/�%P�־�T�kd&��-"��.s�h�'�1(��ˀ��ʨ��/z.t�M�B�/���`�IĴ���~�o��yؔ�����S��-5��4��<cV�ȱ�� �Q~���m��m�<��/~9�︕��M�5%�V���kLO�?j�)��4���T��Y�G��4ǔ0~r%��R/._����A-�1��QJ�K���S���s���a�.�S����+�|��#�M�|�o��$5s�5�W�ք1o|����7 ���Y�;�3z�MԴ��O�1�w^_���~澧����"qu�k0�����x�j~B����2���Z�����;�UR�C�'������=���@Qv��}w�<��=~c�Ok��9�Xk|�Y��u[�Hrd�x
�*ť÷Bg\��ڂݙ���v�Dc�)��xm������n�)"_�å����������s��)��{�t�=`�u��ř*vc�L8���D���f�����]�?x�t'7�V�Ty1tj�{����	B�O�tt������H(*3e�I�6P�s��Tn�QBv��$��`�C+�S��ӄ۬���.
�%A����o����ü;��[ǯ�kN�Ǫa��2�$���&M�a9pD�llPc��5[�R��<>z�)jl��A��g��u�Mu�NL�OO )�繂Ҟ��׿pK�3U�����o?���)=lK�:.�����:��k�z��&a`cUdB1�H䬽�_�A��1�{p�*T�͑K����N>�}�u����Ť{�����N�8��2
&n0ϳ
�y�ʼ�^���n�x$��_QY��/��l����P���<nE�v�C0�$
����6V��'d튆zV�tC�:��S�	%�G����B�Me�Ǖ��Z'Z;lD4���<jz��l�ܑ0�Q�=�DE����D���}	X�_�q�v��9tvck�E��J�C�^����-�D��K�1]��;pg��ed<�
bٸRܧϝI�\�"o�en�`����X�����jK	ܞ���( �V�֡U$�FU�I��+
+����,����$���2p��j�!x��;;ei/����la��8�g쫡I�k��y���~��՜@�ے�N#�A���Ƿm�Ya5��W�v�x	��8b�z�Oi���߻зK�5����^� Wk8����Y2�[� �Iȋ�*��r��������/e���z���[�{�ŀqH�U\���Ϥ�I�Β��(����3U\3�q�(�p'���v�Hc��v>�e��Mj���[�W�ߏ�ht*B"�+ji8t/���ECŬ�q��W�9�g;���Z���;���ǆ/pj�ty+�J&H5���l�l�
��0m�!��]�.(),���(C�U�`|��x�R<��pӵӅ�ظ<��|@����K�7�T��u���k���L��9��G�^]�oP���K�J�V��1����*�Y(X�h:0�Ten�,(�s��=���s���'�XO�y�X��Qw����K�i�w��c��~�^<�ӷ�����$��|Ղ���#����r���n��
1
T��N��E�kw�C���������i�ZA�N�T����f �����;]���\����,*�*��%w�gv�� 1%��t�(��S�������6VPg}/!c&�3�nV��_�5���ڕղ9Y�<��s���#�+Nl�&pN]F��4��.1paX��<��稂BF��Vr|"¾`׎�YMB��$j6��c�K��[��)���uu�߬f,)���P�lHY�C�h��`OC��mg⨮�N��at���f����B[�c��a���1ͧϭ,͎t�^�`39�$�џ�:8X����_����l��S���l)��曧��N���6�Irt�Z��hXQ��B��G��e��@[��q�_?'��4{�qr!ƋU�6	��|���\���g��rh�^�Qfx��1���X��L�l@�Z��*��D�P0�H�\��^��X^���m
������՛]N�[T��x�b'J��J��턳��Oγ�����)v2d�.F>Ugx�
D���S= E��-v�+�Qγ��b��X5�"�u:��.�W�Ink�2�p�~:)�,�	�����e���(�O���
��2����t����e�^������B�xz�*Jy��t�fR�+dz3������Ƕ.�Aho
bFD�0�Ǥdq)Z6�s3�S?@��R v��-�����^wB��]�Ѣ�p�Df��gbN�C#ЛMOy�F�����[���X'�Q2���S�`F���r�ΜX����3⬜��|�{�Q��znH�B��?����}��p_�{�u�������?��3�H3��~��"��0E�`�\��JlN�X�x�>,���a�C,��z[&��k��g�3�X��ք"Y)G���xf��>��3��6��?��Č����6�ڼP��'a��`3&jNIR�����L�cT�M�~#
���"`�����f]�5���";��u��%����^4�e�>�(@"^�GaU)��Ӊ��s�,@�ӌZׁ�-���Ъ����f{V�_��)XlxV64EB    fa00    2880S�*;9.�b� =ZP�����tAuו��Y��GU4i�b �G!���
�U�s�ר�Pu=*E�8�t���(��f
�|��9�S�c<Ŷ�G�9Kx�a6�F�Ց5�4���IʑZe��j���N��k��k��s۹�gF-��k�+�p:�H}��������f��˅����"n�G1R�9`�b�N)�^�ƭQ؜���CO���G�1v���X�*�`y=rPHc|�S2}�<O��C2u�ѥ�h� U�n
���둲#ȰVe�5kA	���W+:$ �95���7Z_$l���Z�~��]J���o*�o-�Cǆ@_�>���^�R�e���\��J
{Wu�QF.G�4��)i��p���S�ޟ���sI�c�kk����-��-nO�d��n_���De�!k�l���Б������]�Q�$�[���7�Fk���a8��ЁT>�B��U-ǀ�NiSW'Sg�2��{հ���+�t�]p?�B7��r�O��7Eo�&�Љ��1������P�y4	C�rTKn� f2�u� �	��2��J�����]р���R�*�?�8�>�fr���3=�J�+��������2����E�t����@M��-���z��$�D�V��Ua�us��T������0��,z���)b���
	�DI�1�XC���s~����d�!��H֒␄��4Q��_Z�I,'񗥍ȃ��xI����:�][�S*�`!��\kF��n~2FMa��˰�Ƒv��1u}:�t�2������*|C���	%���MC_�(+�_9>p(F�O�x���k�N>����T�6}Jzp�`^!Լ�E��q>w��e��@���ڊH����F���%~<���s��3{�{����,WT�vc�5��ՀMT䓪��RߍJJ�=ӹhPH�������`Cѝ5��9al�ׇM�y��=�HЗf�#���d9��YssL����N�l!� (���JCc|�i�wMs��
X7l!��2�}����(6�(V�,���V�/+�/2MF�[���+SJ$ʯL��
��m������$WJi^Q��-�ڈ(>]N�@Kr�]�;����T�Z-�M�7 ��h��)�51��R���v���u�<��������<�����Or�L�.W�컍�W۴ƒm��.��ȵ�����@�0��;|��ɳv��*�4�jZ6<�'3��� �[����0/��o(�(���t2�1!��Ȏ6A<��� A��q]��p[��Ѽ:
�1�{�<�����1�&;$53�/:
��R�-l�#��_�C�X��2�A������h�/�\����{�O&��LMf���$���*�O�RŪ��+4fx,�5�5%�Z��"�BW��i��m����j�8�:��U=������ܒ:��pW04�tw�?�A���cG�$� ŀ�T:��<q[�W9�%nh1�3 �M����֦��+�:z�LQ*�r(ع8��(���d�ܳ�|�� LօNu�`�lX��8���q�5p�[����P&y�����9;�6�����q%m����;�N�o1��sY���݁�|��<ܚ�����2#�r���&gt����$7&>R���IHA�H�u����*z:�8�ǉK�����`��{���'�XJ�����h�u7�ANȝ��Z��}���Dxv�.��kg�_�.\�RdD$ܟ�3��w���b�*�4��O�{�@�Ѹ���ܫ�!v���!�5^�F����u��[g0s�t����#T/Rݹ�qG�<���4�h6���TS�����~��с�<�"h-9�5��g��š��!���2 �M��h+�DYȺU��%��aU�H�5�9��{㪄z
x�(9�`�̺���ڗu����q��ۜ���Ծ�TW;sd֙5ٲ�f��0�R��Ɇ��J�Rz��3~�OB�k �]�jR��pz=EQ��J��W��6��I�ǡNPj[�2�NeN?���/ �YBg[w���YO�=�p����Z�Eo��bSP��+G7E=�}1�g)��؅��	P'{�q���#rX�_��Z�A������#3ﺨl����'���Z�����u[�X>���=�36܊���mg�Կ٦oԮ�	@(U���M
}�o� �^�z����[����4	K��q.��'�Ї��	����u��+�!��}eX"�p���o�[�ފ[�s+Ȓ�e�f�����pK�o�\�맩�mE����^1����m�F��t�X��ʌ��\�cTD�f�efp,`�՗EwNk��3�N��� j���j�^io�]C]��P�pp2�*�]�[x,u��)~��S&<���x��-Lg�Σ��6+ƴ���elF'��Ym��ӎX��卋%?.lqd �<s�~�\!�/�\��Ը8��&���'��e�"z'r5=޸D�:��k��S��p-���
��o�!�F�9cbbU�5e��"��%�1s���wMp�O�
l)�;��'V��bD��t���Y�M~���'-t[�Y	���0�H���z}N�\j�a��R�^�v�l
����\���6>�O�P�:�r ��bL
��/�����v�4���<|3Qo�����I�H@b%��E�m��Q�y�s"l��6��q����1�&kLϤ5���v�r���4��a������m�t;���S�t2>�̃�u���ڭ�h�?��[�r%Y<���,�,rCuU�]�0��Id��L�;uWpD�Sź�3�ӛ�v�y��L^�ʢ��Yf`����$�����V��噂�"�!+�e,�u���4�Vc�n�"+�}_Zr�q �Ɓ���Ӛ��z�I��0&MV�ٍ��5�_���z�p�C�L��N��1�ĽX,!��=��+���F[c5v�K}ߙ1 '���$-.~��<Da�?9׍Ƥ*�p1�j�p�� �<Ef��=dE�~��!�;��d�(��s!�\��d��O�Ot�5�i47��dq{����0,JO�?��ZM�/+�)E����m���:3hc�"�4�utw6�]��I� ����b[���r�慐�<��"�OK�aݐ&W:�a90�"���� ��ׅ�����n�B?!��\N�z�@��<�\z���B���H�o�q���.������+�ћ��+�|�.~�廱�q�l�-�p�_�2H��{�|���3dnWX�'�d76�#UjFH��+o���/e�`qZ���/�rjؾ�(^J������w��j-k�M���Hg�W����U��i�uӁ�^�"����wn�TJS� ��:plO+�I����G�6o$�YЉ1y���z@&�\���<X��`
��}WK�6"1�5X���`����� KH���Eo�T��;q���b��Be���zE��K�S^��<�������;��������${ �3��d��𾶾�|G��Sؐ[�A�ȝ�LL�5JA�g�̋8钷�^���`��7�	��>!��F=H)b����t�ߵ�ZgxM�""����-K�z	�/���#���\TU�1gPO�o�X5:�e6�T�/���'�+��|;�J>������̒"�ex':c�+0�Нy�8������A�� 3u�n!������uk�Y	o���E��p��m
�Cv���keF%��H���Y-a�� ѿ"��!�
�"ci/_H�##7�z��8���<���J��Fe�x��q�K�IcN$Ձ�#Z��W��%�-]�k��O/���^�J�b��!�i�S�~��<_�]�ư{�!���*�U�݌��B(ڍ�!�.t�kqi��9���KB(�ש�?F �9��l�����O��b�n�i��~�R�D3q�_����h	��6�z�<��sr�C���v|R���ٙ����o(	Gf8|�R�����r����Md�[=7����fQf�oV�T9:�,i�4+����9���A���Z2�Q����4�8�.m|�kN3]���FR�83	��0ӯ�X0F�pl���M���Ao�������/LQC�۳\�eG	�h�z����� ��U��a�.X����,������L�y���B`�M�_xwF��5��U����5� �d�8�e�^
R���}p�qކol�~71��:��W�v���6���Yc �b�>=�fCEV�~%zÓ�W.~]��e�����OE�Y�Ӈ{�Cn�G��{5}�c�(&�veL�O�K�p��(�c��p�dw���(�n�.!��R�]���YD����3 
;jM�m�|N��7Ѓʅ�#saŷ而�-X1vM��&�.q�}E�nU�7��'O�V�Jĉ�6�6���Q��C�#[O��7&+�-rbZ���+���Kg�������ˉ&�ѱN"�Ya IE�[/*(����7��!Ɵ�(�����x(b~S7X�@�-�_��8��U����o��K���_=���������t�W��[��q����/k��]�0e.���:�������y%(��@N�Dխd(:��s;��}�/�ѡ�����7%��IWx����|6� !9���i:��k���r�1{��]������w�����G+br�.���cځ�l����;�)>�Rj�gb��o?��?sys]ץ7����q���"�q�EX)�:������Φ�m�Ø�N22rP�/J>I���Ũ<�T*��h{#�VwO�\y�-/u�f��
l�5Xb�MzŧO�A3vpKNYx+�6?�S-k��і%�5Z]3�p�"��(rf�9N�JsŖ���~|�Ra� D�>�_���D���Ă�0e�?�������k��'-=',���1}�SB�v!(�ˤ�T�X��W���)� u��ʹ��'-��6w�$6$Q�UT>=��P�V�m��{%�)�]�d-A��� N=z�L�#�~�С$Ń�dDd�js��	(����P��4����86X���Tt�c>+�`I~�nҳ�&����AhMrM�~.w'�:�0�I$���9���n���1�Y|@���S�����D����1u>k�3C���j�R]�ݯ�ŭ�e�[�ڶ=�W\�\d�ppT�v��N�L]��P/R�H������%���w�;�",��D�*�?��r����^��*������� Z�r
�-PS���Y)&·���P����|�%�a��h��3��E(�b��f9VdB+�n�б,{x@pY��N�����j��������h52��Q�r����H<flo�(�
wm��|٣X>����0u
�@�7P�U����>�A6�(_!�5�~��$��%���#�L.���s����9>������I�1��^�?�#���ʷ��N���:\hg��ƹ	f�{����3R�]_#��%,�$�^L�e.T6�~�=�ݵd;�C��H?��A����=��>Tjp��7lF[t(/�Y�[�3�� ?���5Xf�w6_��X�񼅠l?�#=���%��t=	�F(�G����1�d�;Qn�[�,��K4+o��\D���n��IN���*�z��5�# ���ӌ��}���3�¥�}�Q�=���u��:�74��$��.b5{���Hr����>�{r�`j'�b��֪�"7r��؎�����e���N�� ����hf�W���n���s Uq��ܪ�y�,�U�6`�:�̆oq��}O�G8�9�.պs�����ꔄ4�i��4�6Va����:���7a�doގ#u��[b�B�="p&a�l����G:N���L;ua7�a(�q*�9�n�R�̰+.����o������0AI���+��F��� >�����[�P���ij�˷�ː���o�����L8���%�7���]n\\m�k<��,����<��v���5�WvV��[}m��Hz'��k�؋�u��渥�a��C�s&�`��T�@�1�6ix?��ƅ��P�$/����C]ћ'�*�h�ܑ/

�s���VfZ�3g���{)L��t��ȄJb�&*�8;]��ydձA���_���r�d)�$�B�����J5��V殠Z�hOc��z��E˜�~���b.�li�
���xӨUh0����\2@^�=O6ݨLe�Y�>�p��0gyEظ��A����>��$7J��> �vg��ǂio��ՠ��ԓ�JZ���a&B4cn��@�����z��:C��;�۟M.�O���gyP��I�oH�r������Mm��w	�4��:_�^��MKץ���Wh�@D�*w+J6%���f��7L^��hCXmh�w�0��b�A����!����ᣞӋk�,�,�FG��� �o�d��A �'��&�E<�+�W�0r���z(5/�M��[�g��]3#24�vK4��/j�T�H�UK�Z[��g'�i�j膜�_����[G�����YR�eJ����m�e1��2�ғ���~�=[�u��+������s��B� K���ä����P���V���Mmzk�n����	-`ԙ-��8���5���Ƣ�bI w����ܪ���-}Ũ1D����,iO<��5�%����f!��	��Y����l��������T^ٜ���s�[bG���v��Z�%��W��]��� 9fM�\^f�۽`�����-����F�on��>ԍeFZc���B����bW0�Ri�����)[�
�8	��=�Vzh��&�O|����b�o�c�6���2�R�I�F���6ԓ��cnɧ�'2�5�t¶h�4Y��	�Nɵ���jp�Ƶ�8ic�Y�3�d�Sq;�px�~̚����r;� ����|о���+nz��Y���.L�����4�bi�_��Ф+{�53$ U��?����&Цq/
�i�BJau��F,�Eh�����3������T)|�݌�I(�1����6��?c��Ko!Ʋ�.�4��."_� R�e1�	@��,ޥw��fgթ��Bw���C)���=DYڌ�A�l]*�
�'t�?H±��IԤjw��[�:G PjZ��U[���j塓�$)�}.��S�oK����R�����o����}&8�7xڔ��a�.h,s�~[P� H��O�t$D��x��*V�ٞ��#�.�3Ǣ ?�l���n@T���P�O��4���?�����<�˓Ƽ�5XO7�[�01��U(f�	�	���$߬V>p��䉁p;<��U��jʐ@u7kV����~C=t_�}�����1�T�Y�;�5\��m_�"gt��%�(��FP�C�`0"~�Xm�>�8�hdJ��Ǳ��r��̶��	g�hpy�ѓ%1�B8��Z�g����쥄��:t�2Yb�.���U��C��n8(N�GFiq ��r�4��e���R��� a�9��o�i�z�7�����[�ُ-�d,�*�PU5H�@�aM��EL�sA�G0�4���a�eH����\Gq+�m#^#ǁ�a�n��r��lD&*�T�C��ޜX�p"���R��r)��P�> �5P�=�?�#�K8c[*bu�|@?�4���+�7�?s�5��q:!!�XV�X����Fq�7�
�䵝�D	�)�|�eeK�4L}��7�2��܁�w&�ũ�u*��R�ρ��e7jw�΅ �j�����]�մ��7�:|��5�Ȯa02�'�1o�-l�V5(%3��mz���^}t��",%��oQ���w�\xMam��L�wEL)؆�0BAK�kX��k\ϖ�h��wl0��zj,�mA�d-�6�C������J���B����"/��lT��o��F�IY��zҶ?����u�Y���~�l-�O�q�a�A.rb25�Bũ��X%���ҽJ:�y�I򊵓��T,1hcu�c�lkW\/�����/lb�<%B0�Q2�J��(7Z�k�M:;x����B l���[�:���|>zW��
�����ׄ��Gl=�o�ς��pàw��>�c��ҋ�wc��#�:+r]m����c�QϽ��	D=����	����41����1Ăx �-/p�=JFe��d�H�O��"PP����eׄ���)���J�&�'�'�6r��!`VV#�U���t>��0�q� �?��$��SR�;7bn0,EM�dHR]�#bU��Z�
���кA�N��.�7Ҁ���v;`���vspnoeU��Efu��D��@��4�]U�w�Ǥ�[��C⯚�Y@���zե8S����J�J��A7*"�j�OJ+$2��k��QL$!������M���RǗ��~�A�ГH��l}�}7��o7��L���?H-c��B8K���u}`%>"�f��U�� Q٣��AEe������J�XGt�7��J�æ��Ao�fnǻ鍋�4�q^������|�m+fG��ttϓ@||-Ͳ�5�48�	��A�Zw>a��-����p�r�+����u�^2�N��O�ͪ�J��<�B�)��W�Y��0=aS�+A��/T=��'ntd̚�gz��;��s �O����ǟ�>�;
��fW��aK?>朢}5b|j��up�p�~��GLy�mk����`b/>���|��MRD�O�A�Cr�-���DLчWl��߂�Dq�8,� 	���`+�~�a�l��&�-@�M'/�_/�̇'o���e����XY�" 1$�Ok�nOL5����v7ㅀ/�;��MQC�yH��*�O�|Q��\ϢB�}ܕ�e�i:ϼ��N��+6ă$�e! �cD���~�C�]��%8�q�>�~��<,u$I8�ܬ�&�~$�~���S���r_3^�c��$�/�^�s��Xsi��|���&ȣ�<�#%�0`'[/~	B������ud����X�� �,]
�`��3�?)���?�LanӟtV�{CZ�8P���y�C:j�T��7���Zԣ�t1�y��`2�d�ő���s֋&�'�d�L�D|�6��x���1T�[���7+|-�4�z�a����*��]�r/YOW=ő�Z�Y,�%x7��̋>�K���)�*�4N+�35	�FfdۿP����T�v2Ÿ��Y^AԅWO�R��-}H�5���,ߦ|g���2��{5�t��� �w�e�x�쇂oE�d�(�X��^�h$`u�	IN��N���bu�������q� �*����Ѓ�/�S��Ҁ:�!�����#��N�!�)1]̝>c���X�p�-�&=����kɟ�s�Ǒ��u�o�0!��6��6]@��x�kV@�k�e���
!��:l���ͮP�m>�?�:�����	1,�6`��Ci�.��]�:-\y8z��c�[a.�&=�_T�LJߵ�Ɔ�u����C��6���,�;+5%������E�c�t�W�Y�P�e#�R��u�0���{N}�b���~����{����Z�J�n'3�Vӌr�tp������/7����VB��6�!$	��$���rV�]�T&X�����fw͛��_+S�Aɉ���u��|�`jV/�W�f��kr' W��h��L5�@�2�ѥB��۠�j����@�J��b�1�s����0+��߶ɓ ]1�"��xx�cފ�O̭�l��^Z��z��8���_V�_@%����%tv���N|��y��3{4kB��Uz zV���l:��0:���������LV�LT���Q��İOG�����|J�Kqv׳�a\� ��{�I'��p� �*��׵��s-�1Ea��eB�#�4�t���9����7��Ə�\�F{*.�l{r�]�9*��Ď)�>Z���wh���wue�xǧi�M�K�s���t��9�x�m-�j��j�x����tםN �%�!�On/��W]ҢY-�g�y��2�5�:�PS:7^���������Z��N��3���.m�TuYc�L֡��G�#�K����z"�#��d�,���E
��x�7/�O���j���F���!ڎ�C�m.C�ޥ���%e�Y�{{&݂Gm��t'���'Q�2k�l&Y
5�jx �s{���s��6]@�*C"r��6���F��+�#�>t�߄�5����Oj�t��f�cP~�,�0Bh���E�G��@]�%�f3*i*P���[��1��W��<��%jSU���s� �3z���?�}1Ϡ�)nI���=[�{+֖P�z^��5�=��#XlxV64EB    ecaa    22b0�zE0�Q�0�T���a�wp���&�}!�o>���o��+,�j�g����'�f�ߒ�2��19�r[AH�J�I�X�i��[!����*D��0NV1t��9���{�͈\S.�px�eF��f-� n�����9ZBJL�YKS�hu�~=�l��n�+������,<G��2�^��R����<�X�[DɝR@$;���A��������f�m�������&R�����׸���%[rI��C7���|����0g��Iƪ2��>�u�Ӌ�;F���j�`�C)	�޿]�ţ����˪���NO]cf<�~:s�J��碰q�?�ĤL+�ϼ��X.��%��B׭��\+�����v<<��G��}��xf"�&������
�I��E��8�i�:�'d}x���_��������: ��V�Y�] Z��T67t��|�|�O;�ZW���,k�{�E��ѿw��'Cp����v���&Yj&�lÉ���O$�X��"���02���0}�η��EO�ŉN��Sa�Ee� �`F�A�v��6#�&Z�WUVc]F�k�M���0߉Gm�����hB\�w�Z1�|~Yt{��߄��M�����L[t�\�w7�_��ǃ(�D���AW������gD[Cim��P|]3���u�Eu�
f���s9�^8�'�y< p��+��E�y��1�,������6�!�r%
�2�tNNG��RtN�>������I)5���Θ`��$���#y�g��K'h���j8B�ݯ��^���}��lD�^0�4h*�l:���a�����`|Ȯ`%Ie�R�gF�:H�rx�ss���R����@~�,���xyC|���Խ���.��ה��E|`�</Z��Z(6���ɐ=I_+�竁A@�g�k�a>�3�$�O`g�>�a҃O�B�h�f��_/��FIx����3	��u��M�EҶh���"T]e�ҕ0�\��J��xᜩ���yd��4��"��X!fuW�ܵS�(4�Y�?�a��O#��Ny�P
��џGY��,~!@�p+j��ܚp���(�.4���m����j����v�˙���(�Xn�a�r��O�r����5?{'�
��${�<��� ��Gγ�ߙ�b��lg9��#.T��&�Y�ÕO���[}j��;�?D1���n��a�I�v1;ȿ	+9_2�!���VªRq4]rc����m,�D���&�D
V���g�^�wb0\k.�� 㽩̯��sxd��s�V�"��Z7�$+|�=�o�4����=�ʀ��A0��XR���С&7��m���L촂3:?�qݏ�.Vs��'П]f/��lgޖU�k�%f�n/���y��$��(�_������k�1�no�03}�-� d���۶+)D�`�Jd5�ɜ��
h"�I���+��7bFY�[����-����=����(��μyӌ �Ub�b�S�T��p�/Z;=sfX(M'ߪ8bEwad�n�����t+R`(���|�3m�G��W���H4��� �?���n���f��(�f�I� k[eN��2'�Y/�Yc�HI��,e��9}ެ���䱜{��*���C�F��SS����qm��xx���n{Y�>�V�3�O�P,��d_ob~
�s�H�����0	���	 e[��#Pp�;Z/��S�5̵Ԉ���%�TÈz_�>�^�=t�#�J#�D|��#'��/���QI�v���?�;���
>�O�p�<�̴}�k�π������d��_��k�	��&�P?B�tj4�y���֤����49�6T7x%&:��Pu��x�p����)Yz�{X�}�2-/<E��4$Yn��R����E��j��Upiax|"@�S���%���-���u�۫�}7�o���̈́��Y�s��zsa�]'�5F�rq3��TH]KX��d�95uE��͘|�
ʳ
������$n����j���ph��� �����k�@���(象U��͢����j]�v�>e�"˽d���dY��R��S�U�13V<�Np@�Q6��ē}�\�nR_O>��e��lZMJ�(��ן�%��W|j��K��H�y��)�82�C�)8�mi>?	:{k���H�k���8�>�ٜI��cۿPG�ױ���r��-��0b���Q�����m�W-�v3@9H��w�XR����q�;;�k��\c�A�甌-<>�t�ֺ��A�����z��4�r�������HًS3��_0���rnJ������QYt{q1�]?�8�1C��T|{FK�n~΂���=%�<l��y3�Vo����H�ʅ�KVF�H*�][	��ى r���/f�1�ӳ��TV���i���F�jH�I'�OH�|�IH���-W,�����SQ�^����W
v�Օ�����^��%a�6笧���$V��E��I�9+�/*���x8Ε�
AO2MՉ�	�}���}�&�3sEv-��>�؁�Х��v��{k; 7���Vs[��&h��b|v͋�nC]����R�8��(�+�E�J� n���Ĳ�ck��ԑJ�$��^:l��a6��y��k*N}^щ/����ˮ�u��lz+t!r(��K���o�s�S�MѷƤ��Kާ|,x�ة5�oO�2p� ��MB��,�r.�t$A=�D�r�����*~cfQ�=n����LئPf �^h	��? ���|�@��MmAu�Z\��l��q��G�vh&��~%��7y5"�����^�sVb��o�"��&b۳���ͮ�"kA
^�Q}�kh��!����s�(�SV�*`k�E�ˑؔ�Yό���	
��D艽ȏ;(�q1$�ʗ��cV$k�8Kq6�_j��1E�c%�PF�뽳Ō��bn�{2%ş\� 3+&���Lj^��]���A+�`?��yCĐ�j*TB� W��+�$�Wk��\���� p��p�9Y��K@���-�����ێo(o���&(.5�a<�����
/���-zRk�Ƕhɡ�T&f_x�pE�$	6���oSGo���B��:��<&���&G���I���"���i��(oP�R�6��|��@�i����G�`� ��9����\8��&Zf��,�q�2��	�'�P#������U��S�y�Ax�}����'|�H�r�U�\X�=ѣ��~ü����d.�Ó�7��:�j�p�?|+��NgrC�\��j����g~w�
�!}"��J��a6'���p%�Ō�@����
�0篡`׾�h-�5˃�f�@f�"��CQ�Z@��١�+L�!;a�l}ŧK6]� ���5Ǖ��eW�x�$;���v�#�^U�S��b3���dxC9,-�ݪ�ՃtPx� n|J��	�cC\� $�r�	�.�#�K:���/����ۘ��Uwyɓ���:*����Z���RMtof�[���.a{t10��'�sr�� ^�e�b�ɪ�<�L;��3���{ p,�8LB�0��R<U3������l<vԪң/gm4<7I����C�1��:���EN���� ²	s�ƣ.w�(G��je݊���8���h�YV�����R;VK�]#ņ�͉��D��(L�c���Z����rA@z]a��S����<��â�U��G���r����#2���#h_���*��G_��+�0�h~<#),�A�uʮL�/��B����{G���u]yU�!l[0�� �L/�g�����N�����t��cQ��A1v�ǭ%k���d�#H�Ӊp�Ju ���<�a#@���)nm� 6G�n�ء^�m�_@s�^��>ݠP�cξu'�2)�a= ��RO��Nv}�V�Hu_<�֊Ġ�V�O�{c�2_hY*��8��#�ϕ�R��|��H�Q�J�*��R�� �26�4R)��_�j���K,t��u����dݚ����=�xǾM�w|EuK�f���o򹐱z7q(��oO���٤T`2V;��ai��LfϮ_��Kf@U���Tf��g\�_l�?%3	�>Q�%v�T�(p�.����J��8�gD�qW;ื5�U��5V�yVFȢSg%a���� p��y�@���tIyI���m���=���[lS�;�]5�0�^�i�k�t~5��@��l��ۺ�m̗���ӻ ܿ#*��h�����u��1�׉�-R�u��}x%J^��|�<�ۨ=�E�WNږ�7�xG�'J���|��	?U��������"v��_	�
	'�������p�	����3�%io`F�3��c��0���9�;.(c���\ ���si���I���8`uCݖ�~��P�F_�Þ���T�>� +��ѳ@��Z�"�>��2���wk��z rjŢ��||�e��ݿj=*P�b+e���P�՘�;8e.��;��bk�۵��T<g�~�v(PFRU�0��.��O����+�f��´Q�x��N�!��Q�(�^K��cb�i�3�I%�"��a�d+�B��2m_Yb���`�V1њ�n*��1��L:�Z"�ff_�%S�*�%ډWY��Y��w�<�3W��JF6[���b�R��E��g?����ll|��������5��̀؎U�+a�2���=PAGc�m)Ԛ�2/$x3Pw�-��.��ɗ�nS�Q�Gz�KM�[/A�jrW��L����������h3�2�ŌM�P`��R�$#�^灑���u<�b�^=l
~�'J���Z�&3�J�}8݉*��@@Χ�owo$s⅝�4�'��x[=,����Z�#1��.�S�GEV������|AvuM�	|���"b�[Ұ�f��B�ա�ġ��5X���.פ�\�
ӥ1>-�tcc�ɵ�Y�a�_^�xvyT�T�b�۳~)>�/"0Q�B7g��`���i��Zw,�%�G��x(̉]��
��@/b"�����9���
�\�h/A��B����Q����a���L ��#����p�(a�1rd)(�y&�N8?^K)Z�Ukf�� ���qݏ�3gd~I9e��v����G��g����_��䲃�$g$�d8���n���!d$�#V����\�_Xhα�����͞h�{��Jg7JS�x@���35�_L�{��pF��k�>�T������r����F#�:Wm�����������a�l6�S�����z[GK��Һm��~eQ��?�h���.0_f\����k����gL�ܧ=�PO�5~�0%|���Bkh�Njyd5��̝o"C[17�L?�3���7+U�
�@��L��j��S�ߤ��|O�*K�6���Yw+M�#
k[�'��uwHo�%3�|�C{[�^�' ��y�L��%�4J��U�� C�A��m#��y�;�JC�s��Li$�) #<��X7�z��M!H��T����'�٪%�(��㗍y�����2pn�c[�tk5��jZx�HvX����F?z5峑%95S7�Y�5��͠8wD�}3��x#[�K1��0�����`O�:�;��^U�>���U�h��z�ဋ�l�w����w �&0V�c��`ѽ���צ���y�9��%�.��ES*�k�K���s�����u���c-F��'����MA�b v�du`R�=���
R�#����1��_V>�ǀ��$�cl�����̈ZtQ��R��XJڀ���hњ;��n�k��y61l�W����|�t+y��/	G�:kӓ��Ӊ�5�@�Ċ��w�#�5�r�ك�"v�gR��S��V�a�"'��ޭ,+zf� ib}�3����J5�#�v�P�����f̹��C~k� d��9ZPRk�輼�k@� f��3��Z�'� ����	rP܈�O,�?v�\MM�JȡȢ������Q��TR1�
��{G��F�P�Ʀ����+�$b��J�V7f�+�8�'Q��(v ��5��Y�sK�W3�-��?�7aH���e�U���h��_�l��Z0Lf8�[��4[��\��e�� ��g�ޗǬ�D:�g�������AgRz^���ާxK�9n��|�\�>W����1�-�Ƕݶ����x�X��*��\êJ)�ы�'�gMQtp"$�u����8���>�����b��`� �o��#�� ���w��E�mv���͞'ycEl�8X�2�3�\��;jA��:�Y����������]-ݲE�ऄ�uP�BB��M�J�6�P�X5x�����w8L]Ǳ(��,9�~+DV�Ď�6t��E.d�[~%V������7Diq5eY�s;q�֕�oHL��LT�3&�d�/V��aB���6�$�Kc5X��?�ΎJ=�d��̢�M�"�'����9L�گ�@t!tC�裇w{�XB�6�3�G��@0w|X��`�,�������a����?��`?V���������M���Q�#']���K2�x椆��{��pjr�?u�ɵ��m��7��V�I��B�AQ��X�6������*58M)�)棴����-E��\@w�I56�Њ�)H$E`L=F�r�|�)n����b��91�rw4��z����(��t��{$F�����<PՒcI�K�L�m����ť ���t#l�H�~'����"�5͎6�,�Ɛ���H�E_NSELr��<�̥��R�P�o�`ǫp��z�y�9$��~>�
(n��٬D��)��f�֟,�����1�b�CJ~��]�����[x�C����HOV�)}�hR���vm��:��4���W���3/%y�>��|Ol�Vun�0��[�w���+��U��-��+j6K�ď#�F�(	@
�8�h�9����7�D0(���n�	rUٚ��%�\Mzm�ub� +���_~��]������R9�����\N ��P.�z�à�|/d��$�C5.V�'�u;bI��+���c? d]�����߰n"M���z��ɉ�0Z�èj7Wd/��@  �ݘ(צP�kJ.�1F�W&��a��O/7��ô��|���S&?P�{�>32�%���H�
�g��a�%|hJ�UI���<�6F�AX��q��u���r�-�8��7*�<h\���ƺΨ�ˡ����6��/�A���y/yg|0av��"��f�����Y�%�/9����<�7|�P�覩�
��=��n���:�<�����\�?i��Pdճ"n��nzJ��ཆ)����%�\��W�Q#^}0�b	�����O��+~<#,�����v��h]� �s�ύ �G�Eg��X�[�6��2�����H.̂y�*��x0���R��t�i|4 ��..���P�Z�V�E^�����R.���V��	�|���t��9��H	�ī�(3� [2��mߤ���6����WKWأ��Y�p�/B��ڈ�qz�j��#����m��(�dy�T�KH�9b�P`��+/Ǧ�_k;Tb���zБl��\N�k2Ɏ����g-�������ȫ]AZ;�$��I�фd���ׁ���p�P�$�1���i�����*�m�<p[(�=?|&�����-����x|#)|Po��cI�E�Q"�ר�ļ3ط�GH�H<w���]\��dDk����?�aJ�o`����!i�
[����ڪ�N���tpl��E:�`����>�^k��O����Z�]��$��sbz�l
ӛ��0����OM[\�u�^R��Ȼю��!��_�.$	�D�ѳ��Y%�{:Ui�+�_�Gj���P驭Ů�����**#X�>^+ ���u=�Z0�ߩȐڌ���PG���������3�.��
q�b�a�* ���M�=3T��ͩ 戊��$i�M�a*Y���ܡd���p]������<o�UE�r,�|��~��vn���� O�D{�]bv��Љ�0ξ5�4Pտ�a����"�{������c��Sz?I9[K-7���]����u�/f*�C0�p�˅�rdȅ�'c+����kb�r���I/��z	��f�S=�6�8��:R�^���HL�h�=cj�<�Ε ��|�[�TM����Ǘ��; uj4�����m�hS#}J�KD#�������Q���Txk�N�*�"�]_����^[Ⱦ���,��$ A?�fY�q��h�w21�1+�Z�,��ڝpg���x��7��L����',J���t���0#u��s
8>�{fN#�{��&~$�)`fg<}���\y����2�>�Ҽ�B8���Ҷ}����H҇)�4���<��)$�����S���)��Jq�Ef3KE.���	�!ݑ�V\E��P����E�u�O��k�@r,q����z:��r�{}_:�ۊ?L��������歴������2J��v@�P�*N�rۓr�$BO��K�	'��{���?�����/��
,ڬ���ɔ�@ϲ8��^3�q���W/7�>	A�,0pʨd�;�kϠYu���5�Y���q��]�ܑ��v���F �,f2cM��8@�Q�7<�6N$2n�7��?�]�ь¾��=�,��
�Dţ��h���ḙ-����]��� �R�Hc�I�,����z��}Z2s�;�Ʀ�q)�(	�;=��d�--ba��7�Z"X��u�j��N���{��ަ���-��vy	�47�q�E��_c�Po�)9��5KG��iO�.��#��W�'�'��]eP}��A�� ,1!��3�w秞O/}:���