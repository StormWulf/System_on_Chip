XlxV64EB    55d2    12e0���A�),l��P�M��a
+D:I�����=S���%�N[�Q�������n�B�Ϙ�#�����.�O���\2��}�#�YJ��*?Ŵ����Ԡw��
�hCk�D���E�Z(y8��X�β�Lf+)%��Dũ-/1`�C-b�t��@Qf�Sh�9jX��^b�f��{E)�Ü �����*����	��uǿgT��6�rD������9��4��9���Dvd�P�Oz��
��誛~��S[=U:��ġeE[r��`��5��������;{�A�
l�}��Oʄ�u�A���\������CF�1�lE %�tyG���Z=��>��U���=J�P��k*�����������#QHK��s����o�Tvk���/m��3�/���ĳ1Sz2&i+6�[y����M�ƒ�%�&�GJ�<�*fV�ʿ�ӓÛ�'j����{�Z�5�I(���<��_�"ё_A��87���%*��c.m��Џlpޮꕜ��C��6�]��I.0��me����<I��
6F��		�2͟,k���`�c4j������а�oj���,����	D�o��;6~������7r�	nѨ6����`5^����Q��1᝹u��D���Dm�*�����F����b� _�&P���c��{���0�)�w3f��%��ۼ'�I��=���>
?E;��!岽Y*@,Ƴk�9�����~u�3W'G��v!�kN"�P3��Ц�c�蘴���"~�X=�D��ݱ��rNy�;o��M�)rT�U#��p�/îF�D�¹Z�����lr}Ua���5�/����{vJ��Y-�)1F#);�.�����Rd�6J=��-j�`�>����lH�ק���d~�����ْ�$��^W����>��w�=�������#|n�_oll�@;��<G�_/�e�hs!�jm�C��ן�N;	����ر�/e��؍���Lm���a�-��c�i1�ܶ� RZl/���rD� �=�����_���=��N6t|y�Н	3�S�A-��%���a4�w�G�[�@��cI�����=�8JL���,g�d�����r\�B��O�XUcWtd>l��x�t�d,!���*>D(�>������J�5���q�
�h|���4XG�do���.:,���Q�N`�d	�<��@B�%��}�S�
t��'�2�6��B�>*�ݚX�s�L~Kgǡ�3Td�P~L���*dZT�����{�M��|�����~�l��<���]�̙{�>���!�j!�n���^]6×L�j�@���:��e�g;I_Mm��hq���T��2���b�K�*W��9~QW+!~�����V� ��{��=��A@;��˯M�P)�����8�9D·ݼ8�<�@��S2�g�A����p?k������	���BFQ"吾7Qj*a�v�T�W81leO�
��w1��	�t~�y,ᎎ�$���!����="����a�Mx��D�+1Yc��e/b��Pu�56<Z�7C���2�����\�I�^'�Є-����z͠^���'f�E�8ou#�9E�P9k�ݿ���g��Y�+'��oꝼ�fq�	T�]R!�H��V�vzWP�kY[�b��}�)|x+8۱)a������ۖ݌'����Q�I_$Ԙ��pف2:���Ct�����s�7�H����ص��� �OP�����>h�Ы^�J��MEW�P�ʳ�P�	�:��l�L��8;#B�Yĉj8��W�jI���Y~�C�������Z�\��
U��r��Lb]IN�M�x��Ow:UoZ�ʡ4(���E�=���mK��'^�a�RzK�}*���t���`�{�P����~��Tx�QU�̄5ݛ����w����Ѓo�!�µ�5�Ǳ�h$Q�8q�Uy�눳�T����wY����)!���i�S�;�;��S�6�d��)8�����?�+�D�GH9rV��lh�[����p%��13�����O|5��_�(�Th>�M�l�&m�Ӳ)J���Kā�R5<j����J�f����9�ڞx��B:C+���?f8\6{]x�h�i���_�S�����q+Z,�&������g]�RD?!P�=��m~�n,w�G�E�uCYW܏�+��!��`��&g*�5*�r����ik�RM�6=�d���V�W�����.��������{ţ仢��^pE�q�5�a���:D�0�ych�&:��)I*��!l��˘���h9^֜���-�q�����f�{�q�,>9�M0Yqo��Np�j�6��YxGGѡ3�7�8��������s�T0�@
�lB�\�W�QI���k��(�;�w[���y��p�9F�}�<�e�B%� �� dD`5SG���~u崊!n�1X�u�8�ˡ $�" Q��������Oj���5����&*�r=����T���3���?��
��~�.��|e��?�m�`Q Ӹ'fڶ��p�:0ܓ!��(5U�/��ٶe���.�)NU����DRP%|�>�q��j�N6��7SU� ��0�]�����©�P�y�����rnn��`~"|U�A�3��ei���6�����Ƈ�>��G=����h�=�S�N�S�~�#q�S${!�1���Yx�?3�
ۃ�+,>[��5E�����c���z�����*@�ND��m�ҋ��bs\�hB��/ ��
�rT��� =��z�bz`Gs�y���;U�X�h�����}\.���!5�r���a�g�܂{M��s\�nn�t7jB�#�^��h�{T������pcþ6��L3L'���^�V#��^�`W\�%Ak)Zܾ��6�qwФ<�r��eo��U�<]��w1	�1>�y�3ڙ�
8:1!\���,��ҋh��'�y�C�]%9},�b]#�W���&���o�q�4��:@{+�_ͳ}�g	=���٦t��b��#
��eQ/o�M�Q�S��]Eg�k< �n���<�f����v�$�ʁ�&v�^M%_vW��ԧ�RV��
'��ε[u�a���sy;o{t�*`c�x�"G@W-Of{��;|'_1\�F��Pڿ�Ɏ���ŭ�(�:O,[�#-ː�%���}'�]�ܕ*����3[��纫-�ؼם�dua�u�1�ygk��`�3[P�{���y��8�M^��n��b�W�W�ȝ��� 5�f꬀+�u��*V�v	�}�Y9
CX[t�=z�m��e��cD�3� �đ
F��	� rH����B,�EW�A'��Iz4ً��fz(qvBIપ�L��L��=�1�\�7 Xo��u��~U

#�
6��{3d��
�es����8��U��SQ�Z�,D�����+����h�	�?���T��aF�6�&PZ$�� ��5�<'T�#0��dYN������OJ@J���ܟ�ը6t�$����ڱ�;<P�F)Mۢn�����bg�՝�o�l�"F���#*�F�M�6�� ��[����\�L�m27X(���+hpvz��A��e(>�-�{���e)���Y'�Mʜh(zi��V��緇����Vz8��[�%��� Mq�s�.��\�|�5\���zW|ZG�y�h�L�V6�EO�pݐO�e�H�Ɲ������_�'��	'��%�(�[�Ml���{�����t�H[IF���3١n��K��xn��c����¶P��ZѤ��J�7-�8:�2|gȎ�r����SYoVZb��'��9��u�b�,�����Pt�e*��vn��T&,E� ����0Ar�!�Ϲ:�(�Q��	�W�P\��� u9ps8[��Oo��c�*�7�B�u6 ��`�̨�i��2ұ-��Qq�����U���L҆@$�rG�2�x*��C�Fc�UT��ˬ��/J
�V�^���N���ǁ�4J�C^�8�C���<�>5��� ���/�� 6m�v搫|J��������1}�Bf�!�G��np�#~��Y�'��ZR�Om����©���3�quiBY�y�cm�cr��4���6��iJT�N>��=��	�����8���.,�v/
#��y�Ld;ͺ&plɦ���c�����T�:c�=pe+d���MM!��m�N���ܩ����UP�P�95��hO��$� ]�6��R��Ό/��-��h��8/����g��5gw�:��Љ�
�Ub�A�s^r�wʧ�/��!���cE�ݏ��Ĝ��'�ϜInw^]�u�-����f���Ѵ�Vq ���dܖ��5�Zm�A���*��CةY6��L:�4Pe�G��ioN@cj�ն��d%D��p3k4��gcѼH�u3�!$�5��|��e@���F
�9X�&2�ct)�{�;e���2���S��|��kԯ�Q���%��1�۔f�n�IN��\'^7U���1r������'�8*�!h0�cw��/){��Z��3���ejG15����4l�73{�r��p�Z/ƥ�	K�Hd�)#��'(��3St-Wjk�>�\J?��4���|]qoD��LB�5'�641�RG�Vg���!L|�c_�4}�C&h9��>s2�J~-I�֫N�r�6̓H�
:�|1 ��6��?�#i\�HĐ�V(����e�n��O��oE0U�u���*x�/�1�d �%Q�%YR	\��T�qP� �uCױx(	<E%Ό�[&ť��@'��@m����@e�ܨzƩy��#s׶��E�a-ޘ������a��fr�LK�