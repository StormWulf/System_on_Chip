XlxV64EB    153c     7f0�"z��v#��{��"5[�ǎ��i����=o�~8?舑Zi��0�+]s-㮵�%m6&{���0��P�-B+%;��z�� tP��k��RS��}n��徬#l���&�v;Cy�J��T��H'ܟ'�����2Y/ԧ��Y�0�
�����W���@g��,��S�2�"*��`EQȢ\Pq����N�v������5��^Α��QIa��[����w
׆K0gn����\��>ũ�	��3+��w��]R�jLZ���@mw�X��۵��D4b'���?9�j^i˽;iM8��-��NJ���}�I*���S�A�(�)$��ν\Е�J�^RБ�t�F3�� ²_m��a�ங���}I�_W�N���g�?��zw?y�S��}��=�b�̞�:$�&N�;$����Th�{��� ���n�!���T�����u)"�uhZ���"j�Q���a��m�x�|���
1�]1�G��G/�]A�y巺f�n��$kF�C)�羄e�UV�tБ2f���6ԬW+i��O�~	F����O'�h���E�Q�b��Uŵ���Iv�W�nRC��C Q>W�:;�\[��<���a��AN,μăR�D�Jt��j�~J>�[���F��cRBB���,&m�8h��&pm�g�G���BU ���+Y�i1VK���mfa,D���у3ի,�E��&8���`פi������G�"��m��~^��;#�$��|#��N��GԹ�L����v����U�F�O�^Z/"D�M�P�ލ��A�0��?$����2+�4�xkk4����7���d歑��аΆc�A U�*/�"w��E�����7j<-
\��T�i����1��#O�J.� }�3[+�7�}�x���(�0��cL�������;�w��*�[��*���\���]IV��u��~!�msS�Ƨ�q��Wb�ωY�׀;Q;�޸��w��*��}6B
1��]����ss7B�6���V2��������^:ו�<���5��SB_�ÊsY�4�n�бGb8�)���̹eϖ��^Qx��w�R�#NM(���}�Wz��]�)�RF��"���]��*c�L��!
#U:�q��k��Ticv��\����`��QL⇐y��!XOAFGio e3Q!�?�w��9bp�~���\�x}�6̔��F]�h�ms#��rxm�+��h�Pe��,SVkı����VlU��kN`�����r�YH2�P+�lD�
WS"��x]m�W�۸�ŀ�"^H�3�ŠP���f:�Uʒ���ߔ�ûE"Y�uC���, ���������Z[�'��b��I���8=c�w$��>[O*,t1.��<43l}U t:Ix��s]~��S�e��u��������@�x��@&f�\�X��B��¨?r=�t�o��>e��UDw����`=uU�ހ4��:� ��ϋ�#�ٶ�b7ng��*	���Q�8�ck���[)�%=nu=� �rt�������ٔJ���	��S&��3aKA�.���4̠r¨)��2�W)��n�^��Ŷ�X�5;w�;��Y:�������W�nQ�쑶�zH����t�#�<{ ����X̼}�u�$c_��5�E��K{M�ӛtή$�P��69��_a���i�V���9�eL.6Sr�|s����JSIt"�u	���E�u�LDIF�W@��sm�A�������Vn��s=T� oJ����#��X`B�<q���_܋y3W�t�J�9;���=��[��C�}����y���+��]9}��V�7�= �M)��oһk��^"�>\��=��� 5�e��ԭ�Z�n}4DVL�*�Q�������+�>�cA�8L��Q_�
X�O6���h�;u������eD�I�T��y[e]� ��6�ݲ�?�������z���k�anJ�W�
5��^�R��g7�Ie#�K����7u����X��V]��