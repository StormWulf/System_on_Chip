XlxV64EB    1569     850rc�6*�}�0BiB�p#������K�t��U6��}�ܩ�#pz�����ׯ�}G�X^��H��B�i
~��axe�^S��A���Cq 9��(J%'hSNO7C�^;���Ҏ�^o#�R�p�9���'�𥵧��;"�,�)W<`�LSH!����.�[&���@�RQ����m_�nDD(",���R��O�j�����_o�S�A��t�6U�p@�|"��Fϳv
�A����|�g	&����4�Dk� Z��~JjG�&��i&ab��=)�2���{�nbD�9�1,��VƲ9��9��،ld�w�t��(.�9m<�،N���Mȫh�����Q�N�Z��v$����e��~��Я+�yX���=���>��q��Z<9`��M��(ֻmΘ�� r%���5�.��ֵz��a�'�UG9�ӳ��a�usD�j7=�#�$�8���sP*��B_�Pi��Mxk�|"4�āJ�m�6:콓,����l3�mQfm��W|�d�klq���?��II*�~�����-�Q1���p��XPQ��4�я�*�����'��w�fU*z�}�v���9�_��&M�2�;��9�6z&�"�
v7�<m6�s�l.�&gD���������w
��qc8��_s��>�.K��+m����{*���|#�[a��([�/�̰F��980`�CN�ES.6NZ�Zx��$d��\3R�3� C�6��[�]A+�A��R�˩'ކ�/bLNݱ֮[ǚr�c�������)��a�`p�Sd� ȯ����`7w����E8�<Y�9W_H8���B��ĺ��S�D�X�)+̮�I��[������ZF��,Ǜxh峎O�ÛǏhL94�O@z�{e�%���_Zҷ���*Sgn-��W�j�Pk�����_v���x���\j,�z�#$bc� �;��f7�rC/f����&q��� 1W��̋ȭW�>�zj�7�Y���h��O��=-ʜ�d� ���ag���ke�P1��ʒ����/��eT�K�y����p�0�F��l	�CHeg��zڌ\��5�j� VL��PT�Rl�7�s��:3n�0�~�Klh������q�{�� OM��S��I'H��yKC������	GzP>w�b~��4^��kP�SYQ�9��h�?��l� :�d��{!���K�哚���X�۽�m ʰ�hN2byq2n�]��rR;]���%Dsd��#� ��Lɑ����D8��`�H�s�:'f���pىos�iםO�G���t�b)b�%W��2������p�+�G���ș��weֳ<�	fg� 8"uu�$%Mj��m	G
����3��T��U�����N(Z���͂�`
_�ֆ��R��`�r�%�N�6]-Q�P��_h��k5���,��ɞ�&�ՙ���'�f&��m�J$y�2?���],k ���A��>BB�Q��Y������ϔ·�)���˾���1M0翼���h�`��Ƿ;s��#�ԋ�ѱ�q��km�Ghn����*�b�VGJ֞(i���' �Á?��?�u@����ՙT
�:ʇ�elI-�n��i8a`t�2y�"}���\�z]�2�d��Ћt�%?WhE�Q���:��8�T�?>�6m�0.�G1N��%=����	m���L~�X�|<Uu�RH��{j
[,ߨ,�}��O��䋈��Z��
}��y�%8�y6����kQ�h,�z���s�"ߛbq�yeO��t��;���eu�٩':���s(<�A����(�;�d�Cx�6��I�W�h/E7Ң���gl���4R{{f��>k �~C)�α��Z����9��Ĥ�@��]ˉ����B~;_�]�d�uX<%�;mu
8�!� +��i{�3�z���Rj�����2��'�C���@�x� sw��M�P�h�an�u�j������KX�u��6����h�0oK�K�Q+}[��ɓ��s@�w���S�P�M5� �0�W'��u�����i�(��'� O�$��|��Ѐ��؈�=B�,$�Ј��e+�Ja7OFq��)!��q�[