XlxV64EB    1b8e     9e0�;�G�#�yc�!�ܶ���+�mҕWUU ABw��vd��S��>e;��ߴ6)��9�����焠�w�ac����ز���.h2�|�^~F����QK1�8"
q�� �{8<i`�N�.�
�Č� ��:��"%"�w�:#px:��$(��7V�i����{ �+��C���̀�G|����޵��t$S�z%�2s�yP���;b�%�la�����W���5!%���}{���cB���lD^��.-�nj����ׂȢ��+���[a���S^���xMM�[L�	���|�b�$+S3�K0��`~��n?��k�:�,�:��cʤ9}��F��.0�$������D�d�ɽ޵�{դ�����Fqx0�.WǺ�/�+[Y2:.��S�S�LO�˾�kb@y��D��$h���d�C�x�Cu�]��(�'�;��_a�y����Z�fq��C�Ί]�&\��j�]�a�yV��ۇ�3A� �k���SƁ��i�=��ׯ�s��(_	�	��C%f`3ƞ�����&�"�qx���1��>��_����^~���vM���U�q����Эf� �q�0B��u�ߵ���{q�a�h�Jw��wBb}����d���z�>DǁV S6�h�/�?V%�����	���L��ܔ� �P~���S� V�;�����"�h$S�YL@N�!T�ޯ�� ��Hz�g���g�v�C���F�.tǦ��^�����`���KVv��ߥZ��U�^^-��l��/.M ��0_���뾤�2�m�F��7h��C��0����m���f�1�iE��w����b��sǘr@�b\��>Z���h���A�9��G���.�Iʪ�hV�7#E�r
A�+|+���W�T���4�=�.Vw%��*˦:�/bxa�ޮ~w9W'�O��Wu�!�4/��+�(�劵�z�.G�<�3��m�֚<������H����#�y~f��8�u(��}�j]�ͦfIAz�\~�`\Y�E��B��ѿ�(�җC��?���W�� b6�~E�7}��J$����i4�L��K)���m��h�mj@��գZ�6	�[����;�����ߑw9�P��y��H3m�����m��1�[/��ڽ'��"��;��Z� ���(:���Yr��d��ݻc�hh><*wڀ2��tZ�t���VƓh�4������iZV�)��>�F��n>�X��
k-������*�)��K�Z�s���vKc�K;䬬b��.V�x�t܉5���f����-��暿�d�ŗ�D�r��AᲕ���V(��&!7߆j)��`xS~�9�oE�)�AЩ�AN]m�܊/���`���P�s�lʔ���FR�i���ʞݦ�ל-�����81����ĳő���0�/���.=ޏ��ˀ��!�b����&��^�h�m��z�����p%�ʸ����egn�3�BM.�e�qs�0dҜQ�'N��DɆ�<�����F%)(K�R�}yf�(�iW7t=�5���G>aE��$(�:K%���#�}[�*2k �8w�$� �B�W��}�u]X.��N34�˵N�t8��s���E α�$w���dpn�$*�Jb#���g���s�@�y7�:阑��|֣q�!9a�E������n��˒厑z	5ѐ�$�R��ɥCרHI��Q�V��2��غ��9��b�4���{�OgYs�4��
<�����4�����﷩��D0��_O}�V�8��������L���Y:K- #���쁱KJ�u�������2;���
W��QÀJ��$f��[�p݇-0�=	�������0�r��K�v�}�$/�a��Bj^Q��]��S�(`G�%�(Np����Ԗ?%��i��wc�q]��&���E��(�C��#N��Ⱥ�%s�eI�}��Ro�Ǘ`��I?<�A֖N�08ӷ����xgks\�[�<`�y�r��t3Yϊ�m�qb^k����y1�����g�AooJ68,�60��~3��i�n��V��F��0U=�ǜ޾�Nd�<y� n�c J���Q�w�{�㫀�4F3�wy��k���� 1�o:�O=Ɣ�&�YÂ�𾧂�u1����=o$A( ԁ�E�`�hSP�{)v�}\;�����i�8���`����p�X
�d%<d@�yf��@}��V�ޒU��"+���_�P���Zr��k�$p7J��B��,�<��j�pOy1�5��C��c]�_�O�+MV�u$ۤ1��Ͷ/:`&H���6s���d����{Yw��J�$�|q �풡���7n��rn�GAi�RwK���C�Z� @5���p�Y ���1�
�Yf�nr�`�Dl��@��8�������?��o��@'�+@�<�'���c����x)��9.��G'�C�r�ُDcСڿ���F���v�J��9��U9 ���=Fz6�=�]ڙ��r��:RH{¹�R�]C"