XlxV64EB    b8a8    2370�q�����h8]Z�nYG�W�	�d,9��Sr�+5��űS���@������UhE�|���ZO�;a�#��B�înO�_Uuu�����΃��'��Zy��*�p�M�G~���q��A����tc���~����kۭ�����_�ҫ�O0�ٹำ��ȉ� �b�(��%���m�L	��~���-���Lj���e���dWF�s��N���}�?��r�#�kp>�~t�r��S$+�* �g��(&��W�������G�s��7�0P7�#<^�����&,@���f�5��ub���0(s�jj-��YHΨ�K�7�8��0�Uv%M���b-?��t��rݟ4�#2?��=s>ɗ���l���-I��͒	~�*>��u-�"8D�Ȫ���À���K2L�a�h�� vڟrS���i����m�ʆj�Fc�[aFK,L�7�ׂ��K�C�e`d=��uf����z|;#/�p�s�Nk���,W��i$y"�#���	T�� �ߍv�-+��=n��䪾�UMخ3[e����Q��u}�9�@�#�>!ʡ�7:�V�p��	xƱ;��k3}��Tzs�|Z��}n[���"�P��^�7�^�&�� C�Wè�^`�:!���+�U�g���1@y�?�<��8f�����X9�!{J�L,#'�M�d�q��{�kgNp�k%���}��BH@%���&��&�5��� �:�7���|YTJz3�����̩�H�����!������$�\SMwB1�L���#*1g�c?D�N���akh�U��6е��Z�i�`JO�Н�tBEF�D0ji �Uf[Uז�P����
��i"M
?�9��Z�#�Ӝ�?�5��K�m��"� �uWT+u�N����a��r�~y�ׁؘ�]�M���//�]��P���.6�59��(@�+�^R��c��!���~�_F�����X�@�q�c�/���`����G�p�������u2t��91�j�節1]تߪ��,0�=ZX&��F<Jdnn�>qB�i�p,mR�~Ͷ4�)D՟�	��6Q�����j���$;sa�W~�-lj!��Q��� Ԃ>�Q?O���j;�Or֩N�̇��vK������S	��/�(9�)uD?TK���0�N:q5�+�ɖh�kq��;�0 �X��OiO��Xo��)��n�A5���m����R��kKs,#�@L	:~U9|�����B�ݷ�E�+���H��j@�{�������8gz,�ŭ�͛��L��.Oȫx�����.���Qb�^�T
����@�H����D�ӘdϤK�������Ol�߆�g�%̋v�JI͍��u�_��uXXF�@6����6�V$��"���M598�4=Z�S�P��lAi�[�8�bi�Iw6S�R������}��i��R��S�~�p�-$�9*܀#�8������g�g�Z�3z��s��k��@mvNٙ�`|���8,`�fy�����IO
�Ժw�uq�����4÷�E�y�����8S�^o�q�`U�9�$�C
z���<�]��L�fi.�����˕/Ԑ�3Rj�����B���1��҂H鯀r,��%���!�A ��a���o�Pw/���Q[�I��&`(����1V/A��J6!+|n�Wϰ��������1�|��;*4��(<��2��q�M�d��i����	�'��)��F,}�{i2 e�۵�q�eD�幜�
.�{V�`�*�S��`��{�\
�� �S��(�)�EQ�k�Fb����w*��d��Ӊ�6Q���^�!vezZxTeo�`�S�I}�E�$��ׯ3��99\�{3!��!�&O�>M���,6�căӣ"��91�Y�U U0�|]�Ք�1��i�e{=Ѹ����o��(K�4-~��2�:��g����{�)�]�X}��ëR�彤��.��%�x-Jۅ5	SK8V솽Hm�6�����d���~{�F~}��5���6�4Zb���
f��Q�➓�J����T��ի�-a}�KF�}����7f羮A�{S6�?�"�M�4)N�bQ�����y��V�ԛ�b pB.�.'~%K��O�g�1�Ft7|�td���4�Gfb�Er��O5	�,�h� ��� F1�̱�7��5���V�]=�͙�Kv�|���)��ٕ�j��͑o��B�UogD� �QO3�zs0��{c���fؗ�ݑ�徥�ԙ{BXv0S˄�mN�V�Ъ��X�*���f���	��N�?�$z���������w�Z���D�) Vm}V���Ƽ.�ɴ�����xo�n����݌�FӁ��Fkܠ7w�?�BU$X{*�[��(�����7jf�kZ��($�Y����o V�Sc�H7�8i#��|��:J�����3�ϧ��g	�uaz`%�^աw1��g�B�Z���^<,��D��S�x���`��I½����o*o���W�JK ���Ѿ�����Г�
��j�WLc���D�y��]�3�(B�6SgR�!=b�ru�j����M:�e���zS��w��l���=9c��<	�������z��s7�Zٙ�"�|��
>��p�k0K��a],r�,��Cj�e*=ޅ�V�3������i����vUs~��6�3
tf���Hjy�<2]!��֬#�
����?�O���n�`���-ᆺo�0a��˃*/k��fc��K�Ǡ�}#�Q`����H��`� ���B*u�/r��E�Ϝ;Mbs���i����\���n&�����No@^��=�(n<��~��x��ŖQJ"/��Y�
�u��*���}�/ T\گ�Cl,SPjԞ��(S-�ca�q���E^�F��(7� /о�,��~�� ����7l͓��ʔ���p�^��g�5�S>�K}�߇�az�s�9�I �{�F����(E"R�����i����������g�?�
�k��$����x�ȋ�IA��5��.�tUK�s}���A;*"v>Yo���H������7+��H ̙`���G�"Q����1���MB7��@��}�'	ݵ]��X3Ω��B-FԮ��z:����h�yIh ��uo��V���;�D��K�/^g�	�Nϭs��s/R	��́�(��&h�d��s���n4p��{�q��y�"4���pY�8.�� B�)4�pԱ����)�*d�ˇ�~��!�x+Q��E�8&�.{����bQۣP?�0�b���G)ĵjr3+�G>�J���1���Y�"k���=��$�t�wm����b��5�SI(�Y�!7�EBػ�!�����Lu�a������_����[,�@Vrz�Ŗ7Ѫ�2{��x3�wBp�C𠍒t+�߰'6'@ ���O���F�������'	�O��t�B}���Y,�%מ�[rab���5J�[s=�8���"���.�xѾ��-�-C���l���r��Bo�����QNT|�| r�`Ĥ�X��M�*LV�:>�O"��u�\ݕ�y!檫��р�`vfwT"'^�*c5b�x7#AmwXk�:�Bш��k�Y�5���*�߭��!��_���F��PJ��vv[+���4�g�얉�n������s�El��m�wG�
�m2�bc�Y٘b����#8z�'іN�v����h��O�ho�q��q�:��N9_�M�ΉD�c��	M���N��И����=���$��g�!�R��h������ۧ�u��8��t�4�b��4oPE/���)�e�ڰO�H%..�P -��8P�Y�]hĹ��\A��;��&S��da�b���/Zp����-���\�b�
9Wڒ���c��y�J���!S �
����0���#�ؿ�&�>��<{W��DV@�c��v�E�|�]�1�#�ז�i-��.f$����t�{D���Ҭ���'�YO�0�e��c�LO&1]&[��k|����7������S��=�2Ӣf�hv����h2���͙�m��=���0�_���j��J#��FZ8��pE�6X!8��t�M*֚�s����t32���]!ۢ�X#6��
(�����(�x�g�B))�ĵ�[���g jQ�~=@(3�xW�Kܚ(��O�&R���<	ro��k8!P����W���ٯ�5.�7V+�+Eb�gxm>���p�@��p�ƈ�,�4�.�3�<n�絀9�����7W����
��֊�TI^Lx��E�,O��v�e$����F2�ib�š�f@������zF���JPh�ZJ�_or��m_��Jd������tp`͔�\dO���t�1$�� �hW���J��+�g_[�}଼ �!ދJA����͸��/-��؏ꃿ�M���u
�����K�e���R��D۫D��G6�SGV��HƼ���R�Uص2���0����PP�.�C}�Ϛ�J@������E��W߅Ok����oRmj�8��:<� �Z(�H����7�����5�e��	��\?���|���"K΍�;hr��ڐ5[̵�S�#���n�P��J+Pn,��$��ZC��HUv4�߯����b+h��S{Hͦ,^�ʪ��M�yK<u�O$�y�!�f��p��:��D+0��e�����g��J�����JT��ᴩ+Va�#M�/��`{��u nS���}�##��+_�Q�Ws<>���sR�� )Ȍ��
\7[�S3�H�?!��T�:� F�����EN|�ci/��.��G�m8�P=�t%Ár��Eo=48��RTH�������1�éa��{�O�`��4#�ۘ5|��K���Nq�Nʙ��:��)���=���"Y�l�y������Ҕ�<Cz1�Sɐŝ!�-%S�a�UU�T���y�0Qvh�ö�`��L�x��C�,����"��l�J���8>��8�m)3H�XpX{�[_ɒvk�|�y
A�o�s5K�X�����v�������VM��is��5�X�ᤧ+7;Ε��f��ֵ�c����bÙљ#�,u���"�G�>4��λy��U�����G��p]P�?HrT5�;�hxP���%�MzT���뮞Лc'�4��H�hX���l�5oT"e.�
e��X�D�����GDk�a(�W�8��o�#6H70F{��]͖�ǃ3F�g��j:��LyD��ųW�'tۭ���gOӒ����c$P-�����S�$X���=+�w��T&z���3��љ�	xPO���|>���wYl�cW�.��k�,�4��0��g�7�p��� �6��Ͼ�O���cm�=�;�*��hq֩��K+�x��f���o�q�D?�y�o��!���������+ߌ�2r�さk���`�S��,A��Nf���Ӈ8��At~����Q�N��u�c�d�������n��u�߫@n.�mȀ�-ݨ��n�MD�<�k)"����@����rp��;%���n]�x*b�ޢ�`ה��ڷz	LĿ�|�V�����@i��i��@M\��O��7:���*��ѝ_a8�s0����Em	h�#�߽:b�H\sv�nXo���Ķ8���Vh]W��} �.�zP�p�;�7��
8�CFa�/�J���{����ẘ�Yw���z����U�u��>4�����QTo��ݬ�t�����	�$U�`欀�@<OƪtI��ݺ5�X	����[/%����g�\k�c�e1I����o>�q��W%���gT�����C��_����9[�^�M�L�@S����3g�;B�B�u%?�M){�	��wL����zk��b��T�����Z���a3KtYwʯ˙���e���e:5�R1���I��rҒ������|�ZU���@L�+:^��bX,a����Ujp/+�^��c  -�Q��P��;|?@
�C�M�G(���"7�1����Yӱ6�3�g�e�3N2�7����c��B�r}��h�t�J�iKݣ��Ѣ���d>��"AZ�����<K4�V�wd@���s᧧���f�%����ǡ*J�$}����J$�}����R��26�����"��6 �
�ཀྵ�/����0`�9���_�2��&�Q���%�γ��0pD��u1�a��S�ga�?�p< ���q�D�������@[rtxI�}��vw�\!Y!�a�
�7Ι�X���V��qC�0OW�v�EfQ�o����_KB�Ao����]��G��A��g���Ad~�jI����si ���
�7o�@P���d@2�\�i:)��҃v_-���<���(E��*��p�q�!ʾ-��R6n���Q��`�"����~B��u�E�<="���{��F�:���O��W���OW��!�J�UE����هvGZ�Ӣ�<��uY����@����خ��!J�k-4L��,^�f�3�o�m��C��¼ň(��c���R��p�Yowᵘϼ�`����+U5ɼѸ�f�+��e5v��{4�{	a�e����~ɸ�*Ҩ��|N��d��O�P�R1 *E
4b�<�Y
��"��1�@�
�e\�1�?
�KM. 5���6�u��H������H��_z����	�b��l?-e�M%�J�o��ϔⵈ�b�S{}�+�<rx�E
����uٙ���"��=)��$�t5���w��,��R�PU��̗��I�8~���p���N�,�SCq��Y�N�n��f'g��R\��X[�'{�e	.H����a�X����n
>�^#`s P�Ϧ?��Y�e�1gG� $�X�Zz�h�P�f�B��&��-~i�>/ˍ���L�3Ϻt��G�F/]�SKH�dvwG:ż]��Rl��{�6hf�^D�qLk0ҕIE���>I4�r4؊�P�t��M�è�L�����ݻ�/����L�����)Ui#�����I�+J˯ek�ߠ`֗V�5$^(ĸ&�^B�W�52�
�S������+N�沇tDBf����47�rSL�ϩH�F>��ͩrE�>��X�)����[�̫�H�]K�,�o�����`�m��j�5���h�$u���_(�S���"mm�V>pa��a2K�9p~�yW>rA#(ɳ��-?`����a"�1CJ�Jr�;�h*��[����'F��Ej�������"���B�ש:�|�b��TO�Z�������%����NB�3�V8R�
�`�]T-���.�VU��X�A�ފH0��m���bkMRm8�0DHc"ȠG���$.�T�I=d{M�7���r�yw���N熬�w[��_���76��mQ��׽� I����# D��2�. A���b�����Gs ��$H᧼?ҧ`�����#='�%,��f��4/;�>���v3��6�%xi)p3b���I�˯���r��b�}S,p4'�Ա�Λ�@\�ŗ���1F�98�����Z�������TP'd�✔h��'�W}lI��8���4E7/�0���ܕ�	������f��~��K�qO`E>X���o���J䁺�8�y�^��Y�7��qmPh+���/���U&�z@���Z��Z���ʦ}|�� @XQ4VBk��N���<�Z0ܷ����!��_^Av�M�1���q��?P��T��F�;v�\=�=��ٌ�MGx��L��6�0J��?�h�V�����6&��q��:���5��z�V�˒\��"�:}k�s�m8Ōa�����<Hl=����h|�X�`�d�R�G��"�"�º�	v�Ϊ[(�˓��'���We�ѡ���/�'��%U�IH�,S+�1�7N�_8DL>qs�(#�䘵n�e��ۑ�*ǱИ��sKw&M�p���&7V������s�r�km���N 8,xH(����dx1㿺�'Q��	�s����Nb��~�/e��cA��LjG��,z���`�t0Z���>@*�AhlhЧQ2Ca3��*�����6��|�S��Q����(n0u�����B�w0����jL���l���b}e��-w��oU|7ZTa(qSs\�3���On��Z���q��Ԃ��c���u`�kvm��%g%��;�@RR�d�ŉ����v"�oK�f�B(�	=�r�K���9_R�ǚ��[Ή#�n9�1ʍ�XL�Ȭ�[���b5���N�v���K�Q`,Ѭ�"=���&~m������ʆ)��V~���t�9q(��b����u̅�2�����K��w��r'UdJ�.�t�Y�ݸ6�r_�W�0j������6��U����{�}����Mm~�-�8�mD�r좚'�ڜF��'A�������")�����K3w>21b�w���_��I,���L�����^�:��4_����sL���M��.\�I|<�Ң7治G�f��7?~Ii�~6�e��@5�Z�F*�l��O�L��:�Y���&4aٳB
3��	rUc%�ur�#�²%e��wX��W�� �q��5g��7�pD�x�r)��\�h�|ȅ<��?�l/��+(=Z�$�}u�	�M�n�D����;��܈�-Ȋ
c�~a�.w��*�U�H[�)�
��»���Oϸ���s��ƍ��T�X���j��J`G�SOW[�Z^��3���x�n�IR����]����'|�eW�B��*�?ڵ�Lm��<�W-5ōӎ�\�r�q���CG㐿��c{q�z��|,?�_��d��W����OgJ?�R�$B�`�$�V��t����՛�b3f@簏V���ZY��2У>�'��*aq9������9��J�D[G�L㹵�j��6��Rp�f�i<y����u�8�9�� gt�TM�b!����d�����K%����_l��dyl>Ϋ�>�Y-�$��� �(���k�3�m�қ�Bڑ�Lrݖ�F�