XlxV64EB    249d     c60UJ�?_��X�Գg&J<�w�+�[�T�ٰ�������L���?hߍ~Cd��xÑ.�6��A������� , �����( :e/W��|�&��	09Ia���n&+?R��m�!��N+*��������I����ĵ�%wI��mBlml
�F�К(N�<l����	$���Y�v�T�V]�}]��~�7)�0y�j�_x���w|`��v�u��*��p%��TB�V�T���b�û���㛒�oM���w�����L�}M7�\M�N��+.��.2َ��ȿ��5maxVj�m�����A��\�ͥ�$����ۘ�w>q���ڵǍ������E�����0[�ٶ
�8t(�[X�04foP�gܑ&��Zb58��!~�|Y��t�(��pVČR
h��"��:�{3oIu%�k+�D`��E-���yZ�r3�%��b�<㢯���&�:�A�fV��	4���um���ﻂ��ty���|�����2>���t�_��2�4�UlPi�Vf��_��u?���{�5ݎ�p� a���X3^�d��Hϖ���T���]C�@��O��ge�S	ԅ�����xb6�S �h�P���U��b���k`���Hj%�F��w�8é�c���'���W�2�N���l4 �*�`˙M�G�y���^L�MLK��;��$��M��..Q�T�L���!o݉�c�|�7�D 5��`2L���k��cH��Q���B+K!�Y1~����ҿh?��O2��G.���2۝��P��Ͽ��Q<��|0R3�S���x&����̖�	���<)�嫵�t�%���&4�8��s�f�П_��}A	��S�WW���E�������{h�*��[����\--�o��ͭ��hg^'������3�}�p�K���F��^A��+��4^�]�O��&�"9e�-���r��?��w)�;���ey)�A��� �^.?}��NM���P%!��>œ}Y�� rF��J��䰝f��-Tڋ�K6�>�9Ӌ4W?i��2�u�Lc��Q~�ܼ���IS�Br�*�!P�,���ِ��7#OѰ�}�j���a��k7=^�݋�?	
���7f���:���gɩ����L¸
���ܱ>�!�G�$�w�#����Hy�\h��1+m���īnb�:Ʌ�I��)R֯�=� ����N�g7����e�}T��H*��'1;姾�g,�v��\@�Z�*#Z�U0M)���El[�E7��m�3-h[�]�؊=��Yz��3 b���[9V!�҈q��֍�-�P�\�d��H���ݹ{�8��E�ԥ�����k�Y�����<l놶{{���y5�۽ݫHR.;��3!�C��X���5���TC�̢���>7,9���6�3�Y�f��}RF�j�f��s�:7���={]��.Y�� ���h<7M<�[���l�M�*�"�^I�M�i��3$O�@���"g�
��-�~��0�f�t��Ԋ'�&��4��-3�}j"�y1��f۸5Jk�7���V�b�P8�ɦ�b�.Z���ԗ]T@�������\�����߬[/(x�`%C�c�3H�Zj��<�s���>/�0Oܵo�1���RS	^ùk�aK��3�y���D4������}��C?ė������JLt�%Y�p�/8>Ee��M���A̕�Ug���3hm�&�5r	�j G��������k`B*��;��B� F�ekM�_2��^1�H�V�wLwۇ� $-���5��:C���;��
ϡ�'�[d��з�U��R���D�����/�f����_��Ħ��b�4�78�$�>a1��'���ojvZ:PH'L���49ǽq"ä٧�C��P;�)\�����ץC���=�RS�K+�3�p׍�H��8f�s��-���|_�P���@�9��j���2��4/l���������=�^ujJD�FD-;�+_/Z���B)x�U슛�X(���EpBP���x��̱׬@|�>Y��.�0-\� 6'�3�9�,��|�uԻ&�{��K�v��(4I�B�֐o���^�"�#XV3�M�"��L
"�U�y]��R����ZAJyF�]+��4m��I��b͡h�ג�>m�c�9����aXR����}��Ip���[��m�-��4}p����X�脣E���k?�^�_t��5HW��j-�[b=� H���
á�Db��9�
��(�c"_3����e�_[]U��FL��^UU�u�V7��ъ4"E���J��,ZMN����G콶[��06��u��5	�V뀷�����ו��Q�����+~-S7J{�!��ߤF��c��Mk��b�j�
cy��P���d�u27�N������U�B3WP-�o2��W�5T*п��40='�U�Y�E��b� �һD?659��D�$n4�r��1�O��9Nե��_�s*�f�Q;�4zЭ��O��Z?�����4�Wmu��{VZ��ҡ�������ͽ��4��o.+.��M�o�%љI�87 ��(��XRa�|ږ[L S��rHƴ�j�)��|3�I�+�\t�jiV+������v1�%��V�䲮�(�#Af�&Yɬ��
���0�<!�h�'�;�2��@	d�\�ZJ�Oe�y�����bҕ��X� ���FK��+w�>�]8�ü4�T��d}j�9ChM�%�.}���@�b4��g���Pp�R�4�}s�����^��@��������Q��<���O�&�4��V�"\i�"k�jg�pTy�L�p�����\���y�5�ߧ�����5�<���^� )Bl2�;-�b�P�g�3^��ݑa&��!�P�2v�~���K`lݗ&���{��SM&���%� �����,0����2�u�[�.u{��v"=���tQ�Nnj���.D�]�S;��癛��|e|ʚn,����2I�V^Ȝ��o�Njɐ����qT!�x�)����f�P�~R2���̄F�o�HܯKH,9"���c3���Dۺ���,�I\�L�����dcԪ�2����,�~�,AFG���=}�K����Q��