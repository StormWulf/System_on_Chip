XlxV64EB    2706     b70�.U)Qp�iD4pVCu����}Dq:����V��RDaW�°)�\K,dq8n$�*T��N����Yj�/U�z��*�7���2|R�� yԐ%��ZKf9�Z�v���I�{����5P�@6!c���'$lpWmG�i+��?����wy�\m�}��	ؕ͆>e��go�L�͜��m4��P��I�\f��p��`'��I��7�� >�6�@������|N�=��NX5t��W2�~�=@�4��J���ӌ;{4�a?��/��C���Z�]�o����h���~G=��+z`Pb���%��9A8�?	��9�BAz_�쁍䱹�\�0���7��[��	 
 i��͜rV\�6���ԕQ�f:���W��b:>irV1����<��?��^0�>3<�m�/����y��2Ӣ6��
�&)�]�醓�R[� ��9�D�W�Y]�������@i�{���d8��7�>/W�˔������\�(�/��SіW�^a}��3+Zz��)c�~��9� �U���H���Uu�59h��.�v���Q��چ5`�.-�>��M�h�W%���K��ވk��>�I~�����1���q�襨a��Ƴ�r�4�p�}����@˥k�A����Da/k�/��ں�r�	��EQa��[ٺ�F�K/�K<�>aF��K��l�/������0L�&��s'�\F��������0���&�(}�N�̑��WW�"�[r��	�=�$3W�vB4C(�s���>|�rj�ȩ\�R/.8�#����@nz�nE��ڃ�p萠,J��ke�DW�����������}
SE'7�y�J��oD��������RkZ+~dԏ� �y���1.����ͮ���J�:̕�Xh7\�c������Dh%�pq�mP�w�"���t7�{�W�����p1l{�z��6+M���'���S@����{�-�,�{��P#^W��M��In)�������)���KJ�'�"�Uq�6z�1k���22�s��=ۓT�:�{���S���Ɍ�,k9�S�`��җ&(]���PaRљYѕ%88���ͮ&��k*�o�q��q�17��^C���P6�2��Cn $��8/x
��� =�	t]�m}�9V!���#��c���<�е��Q/L��= ��� �U�ˎd%�0�{��K,�H�[D����� q��ֶ�a���|���5�)c���*��!���p0���zQ�'�����Z޻�]�{�_Wґ���B��)���#�ߴn��M�7XQ���f���Gymq��g�Al(i��$�sj{����D��v�g�����ⴛ�pjW���0?
y��R�Ճ�s��B��Q��"`F����c�#� 9r��?���ƞ�f��u�~ݿ�S��`��V��ͦ3���r�{Mܒ���f<\�wD��З"��"O���5J��!�_��Vl�R�T�5� I����'��K��?~��ϋ�"����U�Ў�q%��R�L_�j��ZoNi�ݰE�G�y��aA]Im�����b� N��K�WB��]�Pl|O���½"K,Z�2_�[M�- �����m������ y����9pm��������!�uC�	�	!��Cs?��6��Xz��40���4����5��an�~�'ľ4�0�e�����E�+	K�G��H�
�oW�ڟ���"��R��q��aR���e�WV���T)߃�ӑ`�����ԈrիG�E�Km�bnS�6:8ەU %��1���c�ù���9_��N Q��&�Y�&�����)�J�b6=��`TL�J�d"!�`�KC��(�,���D�X*��돍IA~�����@֫a4���ЈO�u/0t�����'�j�_�!�E����(�3��6
��L3xK�6#��.�]Qc"�� ΈYv�".�T-���$V�p�F/�R�҇MK�Vnժ��ｍw]f�%H�%��kGh�
�N,$V�'Z"c`������̛��e��Fa�����RX�?����z}�ZW5)�`Q�u�MH�כKv�??9�;�S�cQ�K#]�IhmxUZ/�7#>?��\Q�5�����s���tù&:�h/�i,QU��0�yh�qJ�/()-��S�=7f�^�G>�fgU9�̆�9HC�2Z�	Պ������>�H��Lz���GTYءrN��Iܶ�E)ʄ��� �$I��B{= 2*Y5/�"/T�Nm�����f�mW*#�p�ĩ �6��^���V3X��*�fb�Ri٭������3�\�ip��!- �
ߪD\Re��3�WӕK�U᷹k҆Bɹ�V2��icھ��bPs�#҉E���= X<�3�t��^����q��E|���Pq}q�0���8H���~Ϲ��洗���p��wv�rn��A���s�:��:,,y���3?��1)K�G�-�G�f=\4�����Z;E9_H]G܅���<�Zs@�X�N��e�J���w
���!���$^!��ņ4I�����b:�^k/�n�3G<J���x0	���f��G�[3��ͧ��p�ץR���*r��ެ_m��/Iab^@R�Zaf�>9��*�����W�+YM��ɯ�.A,�d"_�6HȭL��<5�R����3�5�t�������GVU���!OB|���ȶ�)ED3������� �����*��g�Ѧ�F:��>��H��v>����GqP�z��snX��:����'��ɩm��8��B�$Y�R��Gmn=�T�~ͯ��q'J����<����mMx�f\�"?(O��%�3�d�2��sI�@+�c,q��]���:���T�X�<����dw ?��-	���