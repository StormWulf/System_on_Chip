XlxV64EB    fa00    2d10���b���=<�l�������>��p�žA��rOE�Hd�o�2S	«�'G������k����![}	*/�j��1�Z��4�u��v��.�9B'\ 7P�g�~=�6��z{��G�C]��\A:�%\��U4���N�����g����#�2�p��^�L?����,S9�Č�����a��,�D.��h�oj"C蓊����}+�L�A%cUW�"�#��'�%@P�� �eL�Z>�=5~���w�� g2b�Y�r�3�?���-�ÜurA��qe����8��@���ifv2ۊ~�׿� �I0����ӿ��z��s�B
(|�~�}#�f_m�F������b� 2VH�!w�.m�$�a0;�3��I �۴��?%)����z�7v�h��o��**RCA��@p4��!�x�_N"5�2c��99����%ʙ��1��O���tö�&4D���~u�s#�1�0j2�����ٌ��	�R���%)c95�'su�7Q��;�礊OYC�tPc.�a^�xJ�6��	�خ���ZW����A�)�K'.ӄz	�H�+K�Y8�A���hP<��7J���E�t�Qf)�D����l*�DI�D<��G#R4���f�ōb���T��� ���X�ԓN�7G�ukx��j��<[bɸz�՟�{�f�.t��&:w�BI��H�4�=��=�r�e�0u������
|5M���`'yORDU�K'�G2�2��=M��LeVO�y� �fyD��{��lrQ蟩 c�(�R��Ι�Ah��$(RiӃ3h�L����E�-@O��|]5^<�H���{�Rj��U�F3��7e��'��
µg�rw(�����E2���yמ��or�����ޟ;��ǥU�V�=�ũ��ڃ�*M�o��@�Y&�@�r]�x�Ŕ����̤h���p@�P��(��y8^_��$WG�^�Y��c�UF�\ C����8��mTU��:��fPD�u�腍f��qu�dH��`���yH/(��9����В��ţ�&�r^�x�M��</-"Dk�c�-�d��cc��^`_Q:��,k�_�_	farue�'�����u뜕�s�MI��G>�����P"�<zQ���K�aӽw^ ���8�FF�+�����~�|s�?���7~Z[}���O��-�/��/�F��-X�.q��orS�(%���3Ŗ@SB��C�7���NYG^��Ty��^�j�!}A���1S��،낁9���3\��*`��'�L)��W`@K�c�.��]�M��S�	�}]'G����7�Vn�*�C���[�]#�6�u^�F`_^ٶ���=��5S�)VHR|�8�5���Jv"��f�	uH���G˯���h��4o�m�#�Xv����9a%+?�!0�[�d׭�8@-�[>#W�W���F���/�ZD��r^':����7�J��Bo�c<��o�0��n>�Zn�I�~�ǔTI�EN��U�R��5_!d�Oe{����d�,���������s!J_h�J���l�i0�Jp�8_�5�;֍{���k�L%�ߛv{�����r1ԩ�������zr4P�V}�B����2��Z#�{��������h ]��ch��ې3ꮶ<�-��2�#t��c�Ao������ D��_^G)\m�,j�N`XSP.�	�3ߙ�ó��ɵʀGQ����ޓ@�{[���5�c��]��Ʒ�8�����i��������K�V��3��߹CO;�J>��մ�4��JWO�PX����@�#��"�nq9s���i�]�Ҿ�;ɤ��D�*p+,��k�Tn�㚌?L-e�:gU�6"z���)s��7�ro������5�րد����#�YCi^�RX��_��4��w%tT�g�G�sIػ;`+s���Ҝ{h!4ݿ_J�����-K*f��p-L(��
q�ũ'�*�]�p�F����:��l��m��[\�÷��p?Y�ۑ�����i�Q�D��҃Zs�SX�$k� 46ݳ���hN#�ۍt�x��Y�[��@wl�țl5�a<�P�T9�Y	���]��呇���؆WM~��Ő�A7a�h��Lw��ta�|2��C��rV��<��&�F��;3W�I��Vkmɴ,����c����j�z00ٰJ�T��~E�@�@�@PҊ��O%
�i�R��a*�<g<?��0�V/��ڭ�"�r)����K	%d��.st@4Ӆ��7���L�,pW"�|�����l#+��kъ~k?Ŕ�<���cBMAH@������A3,Q�/�ʽ{Xe:\�.	�E��-��yJT�
P�s�.<��>cʎqp	������"�겾+��{a|Ę>�0��CG�7-P��������g33���yl��� %�r�Q�{a���F^T��a�����t(��)�˭� ��[N�q�>'/�̵�
���.?�l���Tl!�{Un+Ҷ����3�R���q=	R1)�]�\��=Ä�*e�e�
�M�W���[e�R$v)�щ��m�6�/�!��C ��4}?���+�[�BƟ�ો���w���Ť��	�oU�m�'⭪�zh����n(�
�Y��
��̍�G#`�/�2�ʯ� z�b��)���k<���m�|;�[�1���� �s��R�\*�Z5H��i[�H!�+@[P�hP��Vti��T�����E��x��~�u�
�f!8sd�m���������;4\c�x�Ci��a����)Yy�|T��F����m�f5+�q�E�9�q����X@��~Uw��:~]#x5x�)i>�)ݪu l����c1����@��ʱ�����W� �pr�
�� �Sw�ngʻ%'f���|��%K��]����`����P��Dz���E��C�%������uqzb)t;�ݯB�)}�t�$X�s�v
�C\*��84���2��/mQ�J��lS$E�r�ɿҞ�~�(��5a�ڼdF�D�?�ǝ62T�d���\� 5]�OS[�7�5�Z�q�+�s$�.Y�a7F���L\��>~I���xӨ�\�w���r��kg�[��1w�.V�q��ZR��Cq=8o��'�j��3N�A���/�����W7`e����F�yY���m��Ò��0ῡ�����kV��§�0I��j��`TT��H2��1�׍;�ز�~���_Ho��_ѽ �3A�fq������\"�k׳�g��;��6J�(����(rT�,�̂f�׋��/db�0�"P	Cb'�BX"���~(u����?�Z?M�t�&d�j��+�g��9Kj�G��J	+�B���e򨬲����C&,Y{
��P�*D$,)�����r(+����{*v[��Md��3��>�fU��>�v:+��ĳ�/�K�"Rzv|à���ơ���1ٽ�5A	��]�ٛbE��҇�K���i�h9�!Uvow���8��`��a��p���y4�b�6-�}�*�,���P��($&Lh��8zț7���t�F�ޠ�8<�QN��:l�V��5Q�F�����Z�lM,(�Rf%��L6���"�L�L[��+ }�A��MD��'���b'.P�Rw���K����`��BFRa�]@=w�P�%#�y���mr�-pӳ1�N���k��f�Ep"��Ո���5o���z.�^YΡ���CF�P����tB$��)&�a��?��-R!���+���,����\��.^���5���%H����]�JP�J��$��-��z_�vj�����7�TEx����Z��-���lV ���?�����O���w�M���A�Z%��^�}r�Y	A��Z��>*7nT��h��?�2�-��8���<nP��3�d$�Pk�,d��n�K�a7��꣹��L��Cޝ��g����l�gݯ�2u���Xr-\��u�Ζ!y��F|I)��Q��c���a���cE �My����^f���3x�і��[�g�!�]�[�X�~����1� ������!Z_fe((�t��uc�,Y�&ɘ�f�:Q�w]��?�J�.� ��wG�m���r~p�\ 10z�Y"��6&���>�1q�������ۖ����%����^e�Y���>}��YKj��Z��}Rc|p��Qk�meÉ���FJS Xx���WT�:�w���#%I�Ƈ��#0�#W1N�)�����*���12U�A@��4�7����я���NOz���!{�s������-�?=�ݬ�����-˿u���c�C�sN�E��Gc
��(<y�|mh�W��>�Ѭ�Ӓ縔�f2ꔁ�|�Nv��-�"�?�!=���n�0���9�\ڳy/)�@D&(���O�3��7�x΄�c��L�lم�|��ĔW��}t����b_�
b��u���
f�ʚ�HDh��Twjr�J�/�C��;���7��L�Y9�N�C�3�p�H��{p�%$�"H{k�'d5k��U�%�`��}��Jݢ�����<��Ri�B�P,���!ݖD��eG^,3� ����n�њ�Ƥ[��g�Y�ݎؿ��u����`��cC�7��UQ�l��Ο�)eW_�z��79F�^ʾ��Q��r�����.x�E�_j�:@��w/�C`Na�Σ!�;���K�@����/����G� ��%;+>�f�+x�&'uU�ʈ����Q�b�p���xhR��8����N�T�#{(,ҐI�I�n\�D���j0���'��łi��y�ݬ��!V�e��H�&"=�f:�W?�g2��0���y��c	�kص�?N(�.Gk�LN�esO@��3Y��J�m|�]NOQE��޾��Z�Ob�ro�T�mX!Oe��~\n����q�)/w��&��?�+��"��h"��1ƹ%w4���@��u�dŬ,�ك��e�!�����^�˲n���T��},���:�Ԣt7>�#�wjNU�d��Rd�j�%OR�\4 ����,�$L }�3ٌr-{�F�k6W����)���L�g�u��JX���2�|�S��<aG���6��L!x�E�(k�ԛ�a�MR�3��yj��&�O��Ƃ/S.Z��a5,�1�fގ���:����3�A�5��)3W����˶J�/���b�P]��=Qt�r7'b|���s./"��P���,/$�h-HJ_	z���f��-ߡTpz�|��P[��WNΫ|�V��LU��/Ҳ�����^�	%�`R��*su�FG+l�W �s�X�JRo���� ��,a� ۦ�ǸdR��
�u!-�]Z�9��O�W�b�E}]��i��rB��0�!"�6���/��_��d��;c$�q�w �����S��UJa�$�%2����lan��U��,��|�	P��e~5V ��B���9.�l�^@�e[�i�W^��JCm�h�s��_�z^A�Wk���v8Wi���Gw�Ӷ"�M�)Ƌ���{(.NFt��`����R������:
�l"/��9`�s��c�>��b�-@x��;`��I
��+j{c. �5r��q{(�;��m���w#z�!#����N����Ԙ��f��v���V8qb�^+P�l��f�	���a��+pU	�)BI��w/-�c u��%\�0"LΚ��Ł9�~���w�{Y�sn�2�;M�$��dX*c�	W1k�+��#|��?�OCE�"�_�g��6�!Y���Z�{"��j��Q�֩A���<��6���x���Ε
��j�Ǿ�g�����'RR��L#���b�}Q*����[��ǔˠ5_jE�N��)�;�5�Ij���.ӄP�V(��F��D�)��q��[� G=3L��'��!�JC�^�``)���czY8^:��`�K��fk���65ߗ�C�	Ss�j���(�Yt"-��ATc¡��	g8�f��x1缭(Ɯ��� T�ü����W\ώܾ�B�o��u1�-^F4�#�Qåg��5.�2{�~����LQ+
NY�����#�����#��;�J��R�b4Z�_����`Q��5��Zw	�]^�;�pՙɛӘ�=�Z����-�����B��$����	=&���TZ�&ԴHpV4d�X��ɩt�� �'����31A����+*����>8<�2G��b���	��l����JON�S�=�~a+��@�bi�yi6d���B���$����k�ba��wD�g0U���(�)�X���c���P/����+��~���
�	�pGHw��f%���A�dj^��_X7T�����+�"0�|�xM2�趸c00����r��D'��J|�����A*��=�p�ý*�m}��5�E(�BRu��`fn�_XX)"��s��3��p��Al��T#���q���S��ڔ�5��pޏCyj�(��j�au�<l'�T�p�ܶf�`�]�{E���tv�7JM���c+`$���ʙ'��/�W������M�l���4%Y�X�4��'$����9��(�h���CD2�7ͺ7��S�hl;�j!^v=���
'=���+�̻�:��t�[�r�B�[:�`����}�
"U���kͽ�@v�2���ă)�'L����UAzj�y��� %�}|��e���_�?��A�ftNŘ6d�Y�OJֶ��lсSXҊ���!�u���W1�\�^���k�#.p(h/��x�M���Q@�}�������c�����5�n��q��s
 ��U4CV�X<t 	5����W��]Y\�߫&�h����p�qOd]3���y�]F�w���8��çM۲|�ZN��g�T����?���}�|�����XX��SN��!CeH��A`�7e�B2�_x�A��E���ي_��jx{	]��s���#���/���b�?z�o�����A�tS@��}�oȗ���ô+���Cl+|����@��$�]5/JU~��	ȾF�^x�r]���rhwO�\�~<��P��ŋ�;�G��T�u��?�W6�7��]a�)�kU2� `r�3��Λ��8��{Hę+�L��}c�5���'ϭr�˿:����i԰�q=�48s `��}�ł���AEA��u���6蟄��<��V0��I�N�3�Yǟr��T���{T�P)�����%-@�^a�K5��$[&�R4h���_f٭���b���sG'x�[z�ed��ϒ�^��~�j�@	&L[>7��]��f�eW�5Zł�cHϥ�~Cl�����u�tXD�q�dfXfd�2�|�52��:�^Z���힚j�o7�I]�����j�`j
ɟ��z,�=@O�� x���o��D�]fգH�TwB��$���tp04	�4�C/�gm��/6�~s��j��g����s�q��7�Vn_>�U�в���ez9�5�.ؠ�h��f�A�;�$~/�k���i��cC]�Ԥ$g-�� �/�"bD�P��Gt�����oSl�'a�|P�,��m51�|��{���������(��̚��+��r�L&5�({���v��}��奦V�	h���I3�8J=Sڹ�7s8�fz�y�f;@�~��7��![��z�[p7���Xr�I��J��v�����3�� �<�է..�
��қ�1r�yX��r'M������ 9Z8:^N���0z7��K������갓m�zT'���rT�~�>���
H2 -<)�[g���3���D��0m�%��8jB��tl������$��Y^���K+r
3�>�&�:Ə�U���Z?��T#c���`:�k��q���H�(q���>\ed�s��u�\��j�R��ѯ��@<[�Jw��~��[�~��
9��=�_� ���;�d�e���P��q�?�c	����x�aI��kGJnci*5-�X�
,�f��'(\� �[z��j3��g�E>�����//�&U;Vj�L��{8��i0�KI���� 	�
��AG�7 ��ZW���yoW8J��@�.ή0��z$�,U�j[�J�#��c�~��L�s#L_pR]>��@l K� ``�Ws��{��
�%z�V��OO�{��"|���R|���d�/7y�	�0L1
�`������H>���ε�bX�D�S��$�Έ�K��F��q�Q�3��5�N*Q_��8�L�9(��5۾�?"�Ԇ1���`[f[튐-]��5WГ�1I�P���Kb0`��F��%`_�'E��CvT�?#l{��ҽC�'G�i#סɯG�Z Q�3(5݅�%e���hR��i	��R���s9O)}� #�l�d�	��r��p��$z��S�5G�۞:_�T�WuU��Q�	��h���iv�A�����.D��a�?8T�pE8�S�	k0�_��>�Lɟ���$��傲\�S�_��/�er��=�{�����&,ҥ�L/�2�.�B��]�z�(C����f]�}�2f�@u6�/'�� m{3K�C+*=�N��!�_��l�J���>��b\Ԯ01�!O\3^`~�8�8t�8�7�$��Z�(6c�(Æ�x�(�|�;l���%���0��(��)�,�U�X*�7��1u��Z$�=������)ڷ@�M$��t֍�pORe��z,�^�UO�*B�r��5Y�����O$>��$f��>X��z��kߚ �i�
8O��"���uf0�œ���%s�q`�S-��y��X��5b�y��w�;��H���/�;��}�,�q�I ��&R❗
@�~}C�H�殣���A)a��������K�����A@���/�v�E%�fbz��U��d4c� ���W�*xĭJ��0��×�췃f4���#���̱�������V�ɨ��ȹr��� ��p�%��>6��'y�3._G�����5� [���,{u��n�PqŢ<a�2��I_[��I��j��B6P��5T�0=m��8RA�19�ق���(�;0}m��W}B�k�D
k��R�r�a(_�t�|�/Z���?p9:x]B]'�S�����<����%�:�h=���r{������=�o.� ��/�I�q&���0���P� Qn�	��0��嬽��S�_�c��{K�b��"c�k��$~z��zX�cR�[�E*}��oh���mv��체U�H%�s��w(P�'��+��U��u՜Ҳ�we��=�t���b��@�=!��6zs�'�&NXi���Z�pc��(\���C���}��&L�����s~�-��Q� �ÂZ����OjD�b�n5
pe���Ew��]�'��>¸d��2;������e����<"�?{K�m��<��gLjA�w5y��H�UN��~��i��l2��sB�""�י.ڡ���m��zaK9�� "[3���p4)@gw��3)Hh�r0p��m���O[U�B������Ty��Bⳕ��'���XQb�ǵ�cx|�'��ؤӑ	ڥ�z�*X��L��M�E7*��9�ď���o�����D������S`���6!�v0��)ivP�m�j��uB���^���	̱P�!�U���o�ʞ+m P�C��~�Pe�ϰIǏ�	gO�K�n���m5�~�i"��>t�,j����Tr�BS���0$RW�R���9�-֪�+�7�_�!�N�UK!/��M��|��?
�-*�E�I�F���k�ʎ�ơM�۰��T�4�߼����W�&S8�w���Y���g�ۺ�)j (.iP�\��r�x�j����#��v}�C'/}�m�JJ��(�����������ݦq�s%������K��'"E�H��7��H1����@�8�I�7���N�<2����ZR7Et�Y�ˁ��G3�E�ܷ�"���<#����Y� �d_^R�6nmSۘl�9�!�9��ȁ�X=of9*��.�����DɆTN���؊���,�)��� ID87�7��4���9���d�?(��x�������VeAO��8C�O����G���T�EE�Qf��gY�_�V�B��4���<��٨2}A�W�/����:�����}�g?_�5L 11����l[����܋A:�Q-�u��O�U[�ٗ���;+����� ]��gG ˕߀Z���*a�Fʹ��*-���gk��I�����W�Hs�pu]�ڵQ��I�]�i�>��aT�k������.�¢$���s��z��#��u�x�$`��4��~���������y�)���c��A��FP����}H�^�jѵG-��#rC�<������gH#�V��h;O��MH�򖨰h��y\�e*��۬��Z;q�ރt�X�DsK��5�Z@3�QT�B���f�$L�C��ς��87�1���O�K-*������mL	a��}��b�����U[�#O�Wݾ)��b��|ňY�*�)����I���@�(]B"��L!����� �CsH���fS>�ut��h[$rJ�NiLr��񪢶S�����ɀ�D��9X�T���de����z�e�f�R"s{}4�#���j��;8΄�j�񹐬�Dn� J���t!����>#s�E�1q?K����ѹ�`�om�Y�S��??��b%������l���0�ƽ����ᓴ�r����4�nW�����1Zֺ�}ZYm���X��}��g�	WE�@��h��*�91k�i��<׭��BxG�E���?���x���&*�Tׅ�]�wg���jy�B����i��Ur>�����kn��e�iUz���S����Z�T1!1����B^��Ksbg��ہ=�!�����&�N'���g9/�DcsO�m5Rp��:V����|�-#�.*�x� �#���>�'���#;�ۿ����b���I��7��h��l]8�k�I�g������a�F7�'#[�=+��-��YX"Ҥ?Pڼ�Ľ2x~����"�់���"�F��������On��p�,M̴���� �����V���o\¶h������oϢ�-g �.7I.�U��+H��J�âC��a�s��񦆏���\ύ9��C�	�,��'r>r��3�l(�s��'�r!��$��#`��*��8o��x�8_�[O}ѡ�8�we��Ѕ{��M(=�lh����A�p!ǣBWQ��qp!J���XQ:6��nNsX��iթ#!����[��0��Ra�,]�$���'�i~�6,��������`=�ܿj��<\�8~j;2�߮9��{RP�zF�G����v#��?3p�k�����9vF�uQ5����X#=�X��t|;�XlxV64EB    da95    2270�w6j����0H<�v�X!�K��ҥ#���FX�w*����`q^٭��`{(���ue��8��DE��,�\0����;�s���t	�w�()�v�峹�-v�_/��P����	MUƖ1A^����2HO��>�	�X���B��D�/C��e�މBJ�Tٍ4���>�Xl�*�R-@t)���ʭ`���� �9����̚<�{��������L�>>�P����N�4�!��Ձ0�����x�P%e��M�0�4&t����ȑ9�����g�����v,^J�ZIxo��@7��N�6X��6��B��F�h�N�� ���6�mrM�l���(Z�W~S����=urxIf��f��i,�����Cx�L{k��ƶ�v�L]T|1�E����yP�H����\���[�_31�8),����h�Ph�
�\
�Lf�#1,��ɺY�i��>�Vo��c��o���!_�+	����äu̺M�I��6`�2���{O1s�e�B5Q���C�����7��{��!�k�I���	}�j|`fZ*�X7����t�mO� �������y\��C���=���1wG5Iw���*.Udz���*�l~/e�R�uaK/zJ�I�>ή��
]?)�#�mӉ6�M捰Kry,�*N|=���hNl��8��As|�����̅Q�bn�)�����M�Ƿ�0Ś��?��i���v���~�*m4��z�!�*����m���$L����YTs	`�F�FМ�A���gK%89D;k5(P�~��n����/k:�� �s�DBv�N�}�*�����ל�er]RU�@����y�n y��5�_�&�Z;�|:������B�+p6~���d�ms�Z�VV���G�(w�?Rܗ�)�Om��O���T�k�!V��;����ܻ�i��P�+�5O�|��p�th�N���0a���Rѫ�8x���������:�	}�/�
xM�\�TI=q��s8�\��4�HXFrK�r:KC/J4h&o�{ ��'��ֻ~M����Sl���^;�rɏ���}�4K�o-�_��aM��ah��o��6ɕ��|B�+�둆��Z)��m/���8��(#��~������(���N���Ȕ�<���Ϟ�u���%2��P��sFx�,�""m�y�|���&��f�\�]g>>�֥�MM�>����R�*Ski.�pp����M�ڬ�t�<mLY�?o�j�\����H@�\!!����z�pٗ��Q��B�l���% |��*,���vY;��t��H�4X�l���!zjx��?���C[zq�ϥ�y4�	ޢ_��h�\���̓���@"t���}��[z�Ҋ��wV���Z)�{����Y���ה ��5΋�,�����C}��$:�R4솤'bl��jS?�Z�����2���O�1>�5R��:��[JX��F�u����J�ͱdꐈ?��6��@=��<9��o��Ӛ�K��es��fw�X :U���t~�V*2-@3P�)�@�J��*s2(��b���`��@t��7��T�0v��uA� �;߇g #p~.�}G��8�=��kzP�V$ZDΣ�
�"BڼO�VS�m�B�'�x��YQ��%{�sy���)(��s�wiLw��W�Jc4���ه�+L���H������A6�^!.��j&˯��1���{�\�I�e�����>~JS*(��H��C�>���bk K
��0e$�Í�M�/�G��[�-,�颷K���C5o[��� ��P|�2L�+��\�Ū�H4гQ����!B��{�6�#�_YCV@��k���T������ŗ�IMg�W�@�F�T��e#:�0#/x�W�h���
�����^s��� <A'��HG�F��u�Շg��*�=?�N$��Y�d�v�Bh�S�Ε˃ �{��fx�����5L�~h_����}BUN��D/�^c)����؊;���KD�!�쵝�S���i/�����]>��d���?J?o�3�<t��P�[�t�wH������IV��{�r���S���*O����c��A���=l���#���e��Z8�֎�oz�*jn���Π_�. �?�X�98?h4ֲe�7j7�df ��5ꉳ���1�Lb�X@ɜ3hw)�z�C�q�8���Ak�3�xC�F�B��51�Ns�1tN��?*b��K�U�HE�X.�����J��q:'P�^��t/ݮ�#+��X�>W�Y��\�L2�/;�U���Q��-��dۊ
ý�����%,��A����K{P��w����C�j ���X��SЮ�r[�A��֟F��l������D��@��vI��L#Zη5������j�D�2F>I�IٗmS	Ñ�C&�n�s=v�_7�p���΋�� ��2�������HC�Ҵ�|F���6��I�>F��p�
^v!�lyU�wCp|���`q��a��.��6��cê�6��,�h���HAg.OD�=�vaz�������9��C��t�1$CC$j�y��Que����S������=&���`�"���znWZŋ,�Pú]���ޕ�vz�j���X��P;X4&��m���.�Y	I��).�C0
�KjK�.��4m�W^\�'E���ο�L'I��џwzq����P�� F�ѓqB������E���ݰ{��]c*Z�2�{=H	�vi)�D�<��{Lu�Q��Bq�mbH p�l�R΁+�ik0G%Y�D�U/:9MUQp���Y����{vS,��-�Zw�^�1�j��Ԅ�F��s�H��q+C
�N`V��N��֓�,6�J�n����&��=[��xBm��t�g�ǎ�gO�׃�Tw��H�����b0|�����WG�v����H^ǹC�1�/V�l�ѩ~��gAy�j8��I1��Y~���_d+����R_%�#R|�ەe$���k�I���r�8H�����nz'&���MΝ���S´_.q��nTF�Tܡ|jK��%@���P��G��d(����լ���Y����}�@����YuWS�#�PI۪�h�Jn�hyIu��B���O�I��(C����ʕ�|&B�����o�<���^��م���:���1?,S��On�uڦ���j�[�4G/��$4"���ȕ����D!��H��2�/��:J���5�$���z -:W?�m�@!������?N����ZJ^�z�B4��pO�QO�qx���������۬��|�5�=���R֖��a&��'�ҙ�4(��k,�󙉇���$�%������jZ˥`NĢ�;�)x��>�Y�qb�Ri���즷���w�P��礠�@�骉:Z*Co�Wq���!���KI����Π��;��,�]p���Vr5|���^��LD��l�r|�g5�~^|ρ�g.y����_���Lf��D�2*t�W_b�LP���k�0��bv��L�+�u� X����)b�=՘(����7��H�)㖉�8�/1���y@��R�,-��)ᣄTe-�I�1Mʩ�*C�����H-����|(s܈s]����;-6FCOݦ��@ @}�͇�tk��~�sM��a�H<pE查��9i�IgL�xg�[��ᰧ��� Ţ� ���ɏ����a�칎N�F72t��$|P#����8�ύ��_ك6D�w�6�4W���QlCO6W'ҮJ��F4)8��!���J�./�|4�}�R���t�>0ht����H� &5r�a���5A� �Vl8v�.�=>;��-^� �Y&rAɴ��6�����t��䃭\#@Z��ކ�	D���7@@0p��:[�A�;�z�����+�]~yF*��/��I-���#9�p�����L�k�|+{�.����iǉ�v��i�v��R"L�*���%k��=���s�h�����CL-«f7�.ҽ
�B?؋�<�5���"����H-�>���K�����E�kbO^-�~�/Qv�kt9F��� �U�y��Jݔ�����m����Bh�ꮮ�1���ye��A:�_�J�PC�=#wv��|�rS,�{�I���¤N�Z��
52UF:��ڇhKW_�%	e�������>T�`$��'˾/�D�ZǱA)O�k�Ni��O��E�t �4&_z+���*3��o�J��O��'t�e��|�^�8��Y�PR��o��������RA	�n7�&4�C��V//�B�-�1���@Jk�<O�#��o��|;=��O�:U��N?H�Q�[��`�d
�i۶t랶bIM
Y��70$DC�IX"������<7{�R�Ơ�śOCǇ��f���a����R=���e%�*�CW���a^=,�W��)V��N�[��"Y�nT�uN� �gW�	�K6*��������ՃN�iie�!=��t�.���=9W	�����?TV0��&�?�5)�?S7kN�%�+��@��| ��s��+jk��d��b^���T�&_�C,���E�=͍��ז��(�l���1��iT"O�B�4��	\B�uw���c��.���L*�ͦ7"�ŻدvQ+�}�r,x��[�:�7�@�`$Y�� u���~F�(q��q��p"��ƪ���gw���n|������qSE-/nu!j��޺ҍCT����G�o���W��G�������{��~���h�q6��M>Qi�2���⏛ɥٞU�b�N� �h?sN#��F7>��^���;�I�g���e5�)����N~��(��t��ۛmT_�NZ����:�0��n�_��5���m���ۑ8��"��1&��
��q�����P�3���h������a��j;�7g��i�[�wx���$�%�����@�4a+^�����|$|N�D���a���}��@6yQ�5tO�ᡭ�&��?fz�ے�A(�`>����l�ഒ���t���+�����c���*E�@�]�#�n��F�k0�iq��s7�:/XA�f��z����:��j,��P*shea��A��9e&c$����K�A�.j�����E�4d)�ǔ"�m
:��QÖ!d�a)q�g���E���)��e�*f�.]����k�΄����I����l���)�.�]g,��'d~##!��G������Wrl��q	Bh��d�ˊ�v'�e�4��;��K�i�q{3d���+�^"-�u���U����q� ���O-��U�h�uX�v�B�ޖ�����7\�<�L�H�R]��.@�I~?�`NJ�T�̐M%�|Y��P�����O��^DG���n>�"w��y{C�8���(�e[Īo�����G�W��(8�T��2`�(i���t��:��*c�;e��Y�q���/�RZ�a�5K�e~Z�C�>x3ܒ��q:�Ȁ1�{	�����q����KS�׷a�T�4�qo!Ad3{g.��f-W���Y�W3����)a�*�8��7�|�W3�>1�N�V_����2�ZY����>M��<�.Lķ����o�� �o������bRZ�����y�#�<4����䄣vŨ��p�<Fύ~�>%ǬVf��N3!�l���o����y��Ō��=Ζ+�(5�	���3�D@�m`���Ah��%C+��&�d�@�d|AD$�%�^�v��J�j�]\�����$�1?���Tmp�lܕ�4UΘ�qElO�.�̀��F�}4ʓ��$`��p� ���˨'�vӈ60�.�s��>�^��gq��y���p�Q���.<ң�s������A�ˡ��e�-a��yT�8/]Z)�)�=�;�-��R�8c���1��M���ӕ��J�֪��Bc�@_�����S�H��(�Yl���s�y�%I&҆�ա�����L2�>�dAD����Fu0h�3����K�%�3�� ��ni٠���!3�p�s��Wgη����oZD�˨k��(F��<l�ݽ�-n��d�:I�b!�1�i.�R����t�
V�\LSƷh�Q}�SB��~����R�EgH}�U�m�?�� ����Y��1�li1Ȝ\[����2}:��:�7G�婧�A��p��ʺHQ�ζ���Ek尴6#�ě�I��Oz�s^���kC�NT��đ�2�ᣣ,I��G�2Y�K��Y�< W1E�%}/QNHim�k֙�I��e[3n���`�a}L*+�	]���8���%n��*�q�	%Ԧ�
��n^���VAF�!�g�-��6�f!Q���J�M�7R=`�$��T�=�X{@��ul|a1�G��^��D�J���n�V�>�#B��?���f.>qA��}�Gm�Z��T�/�����#����^��dn
���P����ci���*R|���l@dj�=���A�b�1���AWO`��v��@/�����̔�$�VK���UJ5�
T�q��}8'�0(0�(�������)��(���)�/���RSOr`*��j J��[�-�.�zj�Ku�-9w����˚\�\v%S�"�B��D��I.0Y'�&Tץ�_�o�\�����^��x��/݁�xq�mn��>�8F�$�9�
��9�ݩ/��p��Z�C�9E����`*� ϓx�ܔ��ɱ�5e�)��Et��Z���#�r^J��_e	W��r��C��X�f�v��7�_nX*���1�+P���YXS��>�}�:�a�ڤ�S�u,t����/�-l ��} �Y*��~6��n;�$˞Kܜ��Ȫg���6-Ņ-9g�l�3�9�ʦn{s�5Z��e�XnPՆ���b���1�qWF�j(��/�	��xa�2\g:�,�|�,�&�Z�v�WSn��j��]��ǆ�K�{��<8��k����Eb���Lq� �x��X�Z�0[8�Xϫ�k�����r]0fS�`Y�~?g��Ol1����ے�
�O����0l;PO$nJa��)b$�&��nP��:w?XP�|��:�"u;.��&�(~��2���=�>�Ұ���.Ԉ�C�XO6׋��AxB�i��H��Ƞ�se1_>����ͱmwx\U%O�å�!}�[F:�{�a8{�6�Zdj�#��\�g��y�dh��_����1���.E��/;:V�B�����N'�l6C;e-�y��B�;|�/��"�.P��e%��02�M[�P��;O�
�`Lx6�.�Pܲ�Mj�ŧ�,��{�O��cS�Q9P,E����_59,#�d����^�Y�@�Fu��ݞ�:<�'*�&�����;�����dӖ	d��*�;�أ(��w�E�?虆<���"�]��bY�*�"�t9�sw��g)����LI"�<;�~�cMP�m���|���p���Y�yuf�Uj�K"����@Lӟ�φy���Oi'[�Y+���t��#����?��>hW��Ua�v���l�J��|X�����A����'�]k�Q���<�}�^��z?�@��x��|�q�����K���=��'��Q�6���!{V�z+��vS35
��M���A�)$Ʋ ���@W����ڑ��h ��	%�TA�7��ͬ��P@g�O�������XK0��5y����qP����u�u�{z�dQ3\�N�!&n�~�\"{v��4���$vf��T�vG�G G4&�@.�5,"�n6���E�]��"�j2��dykiAK|��#v����9@Զ�6|��fdγu�"��~�yX�mJ#A�?�Ҍ�|��z`��\C��Ù'Q�Z�_��?f"w�M?�������#��8tS(���W� �W��F�   袑��N"�?o���� � ��gZis��Â��kc�#;�
d/����������m��t��O/qwr�M�w�Zx_�i�������ĀQ��+���WЇ�9S�|=A�eU�����6���V�8�&�]����wu�t :���Q4�ع���$��X�)�*���\!��n�(�D�R׍5�G�:�=C�!nV������4X�-�/�f#�~���!��_�N������������.A������4��H���V��Ǟ�Zc<.��[���2A�oH�Q Q��oծ|B�U�4�k��<��������Wr5@�*�����O��=��V%2�y��e_�ՙB��v ���e���Y�z��k׍�+p�,J�'�_8ǌr4d�_�I��Q�߃����@ªN?�tK�:�3h�؎*xIM�S���	r���h�Z#�4�o-��������,��=$sp���Qv��P�����A���O]O��i��V�N+��4�������{R�%r�=���`�.B�u�
{�~&�M��V���N��
��s��}<���I��en.t0���kK�B���d�,W�gC���5m�լqX�I/����U����!���ѹr8���T`�Hc ���:*�d����%p�`C-�a<o�ɲ-���(�jz�<�3�4�$�o�:��p����[��w���l������
h�M�E;�r/�.���<(���1zȾ܋+v"9��4�\<�Jp��)�� '+�oU�� ���%����P���+