XlxV64EB    5cf7    10c0rϦ�=��|K��Oľ��xwQRT[=�:�L��R�C�������P�#�#f3z�U�ų`�s�^�Ѷ:�)�0>���
V��&tN]"Z@;ɏ-6a=?���/�&,)!K�Z�/�����H&M�~$jO�e� �MR�w���봐^�q�6$H$Ve��M��<��!u(�T������c(�3&yS�Pm�ubfq��%P[��3�pK�MSy,X"t	ں��u�x��S���Y9Ɏ���u�������\+M�4��)�h61:�a�@�t���<��Sk͕����)��`Ĝ��zx�$^���F�d�)_�4�v%Ox=���,��XRkuagr'J��"gck݉���3��eS��w��>uG:{��{��q�JPˏ��05�]t�+%d�C��Y��P�n��9p��ٖ״�=�*(�c��,��eq9^�l��z(|�p�t�,��̑(C�D6�l�k�!B�~��E}�q��w�\��8>�d/����K�q>�%����`��\���EƜ���eR�R���U�ވ����"�C�'��HZB�^�S5ո�����x�o�`������Xx6g�_A����#D��p���Z�����촯vs����C�4�S���|����:<�r
�Y�!g�|���=(�U�z�뭌��YPp���5^ENT[���#3���x�6T�����Tr�pl��A�e�J�)�D�%��6/�6;��q���S<g�c��4���䚃g��l�?��^��oX�m�D ��0l�!�E��c8��u�r�:��ώ�^[��4����(�4pX���>S��>�s��K�:�PJٶ,"��y`V�R��>7VN5�tO��-ig�|��*����΋���I-��!ǥ�<2���ʦ���#����nbG׆�����<+�βo��c�\��O�;i(2U00��5�NHf�s�T��tNz6[���+��*x���ƞ��:Zv`�bl�Y�����c��{A��)����Zè�n��+�B�I����t���Ҩ�o�w���fT3aFv�sGZ���/f��H�N�)!���T�%k|f`)ü�A�e��yF��E*8.��^g��� L&��R�,�_h;�"[�s�F)~A�ˣ��wΫ�܁j���fK�2�FIՓ��]�,Ed�ꯓS�`-��!����|��؆x˱Nr�J�l��*^T�mgֽ�{���L�A���)��3t�'�!���7�(�c)���zw��=ə;��	kL��I�	��%x���	l)�O�@���1�Me���G��F�K�{��B%�+AJ�C��1k��b�PD����a9tN�K�P}y��,�9�����2BY���tw��2j^���=�yw-���6.;�� y�hv���s��l ���z�4\�������E�|�cZQD�B�GG&T�\e�f�-�yʍ��:B5���i���s��Q�#�$ x���v����N!%�dĘ���v��|_��|$\����($W}1--yT��M�'TuMW� ����N�%��Go����9	��^ĉ�v#V*E��|Ƙ�X�q�M$d;:����1"ʀ��ȭ�U�ϋ�?�t|��C����_�7+n��G���d���;�=0|���z�.�����#*l]$�x4������C�w]���ڑ�9��E��v�a�����
{��	�%nz��d��W��U���(7~rc��xq��aJ��tC�z�xu���M�XZ�S_c����:�E��l�ϴx��a�PM~�.����l)	
QE��A~���(�ݶ�n�����ůׁH,�7q�N��@�Z�е�U{�5%c�̦'Ƙ[`�7b���:��J��А_Zղ�o��^��M�o�uvX�Bܧ8t�+/9����H��9P��\4������K���0����/QW�6���/Q�.��	�)�d��=�!8�C]�jo���;�.��E����`/�{��Q��d���O�>��;���z�@�J�lZ�e2��hR�IA����_%X��.��M�A�8��zœ�[hU�]��-����'HJ�Pn.غZ�Z�h��8�C �FV�C��\	+[쪙�ۆz4�H���oY��Pd��RRe�~��@��I���[�2����񘙵���b�Y��g��gF~��?p����W�+g+6)��\��c��_��0p9�'3�f4���,��L�lZ�Eo4�N�h��5�u�4�W�r�9�-6$��0�hK���-�Y��k�y�&=�gի���o~�+K��NyXy��&���+��HE��RhVE7��K>�d�^=Fi��0`TP)�nI5T7��Q95�(���w{��Ƃ7���x^�﨣&^ǥ��X��/���/̋�E��^�\ݸ!��/�4��N�^^��;��9mn]�Ӧ����:��E[3b�I��;����z��:!4�~+��lE>5�����J@�-��ܳ-����_����A���+��_�6=�'��m>�*l��	uc�Ko����
��18Sȟ�PP�U�+��+Xu��I��w0wg�>OR��Í��D�t��׋��T��`��:�z{� Jso��h����${6�#K�i��ͅ�h�uOŻ }4k/c,��	���_$3�Ʀ�_¸צ�go-7�J�F��uK--t{�{ZB�#�U����)�g�-Ϝ�h�sċr��m�2eA��BB, �����o]Kݰe���w!������������W�'��Vt(�m�l��g/CZl�md�T���~�9����R{������ZV�c}�#ȩ�)��v��Z��=zj��H/i(�q�͝�N1��X��b��$��Å�h�.�/�*�uj�MLmJ���"5�3�ak�D�m�ȃ�2 Q������
D���\ـ��u=e"����],K����ZWa�f-�ET�T$U'��]���K���7��F��My�"���A͡�6������\��uF��O�&Lљɞ!v�b�)�LqOh���g����K�J���1��v���pc�}t�R��b��[l���o�T���wDa��j��)�������ru��7H&ऩ�d�=���T�,�7q&��) �tV�$M�^r�#��ȃ��
�Æw���e׌4z�)(,#��]8J�I�.t6M=l�=��\9{�T���&ڒ~��PPy��S��y�z�r�Y�ML��+ҟm�D]87��j4�(��U�
o=@9h4U��-�+�+
�ߺ��{U�|;�݀�˗T����L�������uL����n�I/(<g�ߟ9'���uȚt~>B_c��U�<��_��_�O�>�JM6{2��_^'D7'w
Q�[��(�#�i�:�I砡y;�1����{��Nbpt���#d-D��n�m4�u�V�A��ڃ���JR;���Os���9�p�.���ؤWh��{��@�0q#�P��ȕ�˺պh�����oH(�e��E�<�]KG
���w�C��A,J3��k-�Z�\�����N\݈���$vP%��_�Y4����L)m���u�m����L%0��VnҪ�u�T�V[r��*`f~BG`J��pҍ��yk��,G��K1���A��Q��%���ǜf�u�es�����Y�%��{E>qe��5��l0��(�J�G�A���!V�Pg���N�}�2&d$ĺ�	�R�(>�P�s�Lu�=���G�t~i��ĩ�7�=!�BŜ#��^].es>��U<�X΁���az��\�go�_Q��n= ����E�h�Z�.�����)2�ۥ�ͰӔ�"r���!a�5-�c�� !FoL#$tHQ��?�r�i��	�+��0�����U�R�iȕ�Z��1`K���~�I�ȓ2�Z����4���bǜ�HJ�J150���G&;�|�Fw%RX��myÕY���ZC��b�!��)6��@Ҿ�\ ^���$����W�E��y��J�
��УZn	�~��«!S{$�Xc��	24t�ؿ]_'�����r��CIx��~��U�9 x
L(��_�т��ZP9��@l��*(j�4;ǆ*��!z��>��M஫�M�]*��)I����`�#n<�oqF�
\���5U>�~!K��Ҍ�����0X��XĠ;`���XH=@��_���~SF�}��n#a�k��Wwg���6K6��}d�V8��䟈��g�