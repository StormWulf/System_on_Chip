XlxV64EB    6288    1710��x�ز�Z{����쟚T;s^�y�B�r���(��t� 9�3�V�3�פ.���mnn�!j�fs�e�T�y$MT:-F��i�Z�R�B����`���t���U�r���I�u��%��|�@�'���H[
yXQ�ru%��74���8�%#�P����Id7�C��X�0$-Q ��C��1�K��$R���(+t����rX$۾��G(���>V���x�_��p�7���bR ��5�\�^ץ~���k��i���V�z&I2��,Ny+�x�� ��cH�U��I���9����@��sY5 20��'n�O��Lj�kW�1����	'����5I:{1�~=�')��5aV����᪄Da >%�"�hz�B�y�����Eo�IUψ�q�B�.^�Qv��,+T�,O��ƌ�X؈z>ں����N/!ug[o�R�"�3��du�yg�#~<���Iley8����|�|��Y�_)�iRNp{~����|�hm�|�5�%����CT�;��4̝ʘ��n��9�_xO�D6{P+���7l�ڧ������Ud�$�յ���(�M]�]��ƶ8�9�t�q}l�n�+��`�:�tW?r)�~��n��=+_� )3n�@!�!6��}�J��9�5הo\@�3�[�*-��b��Ք_ ����җ�����7e�ۖ~+��շU޾���\t�m���(����k�EDn��y��ifǜG�+ 	�z�ŀ��'��&U�n�x��G��&2�ߐ�|"&@�i�[�� ��8X�߻s�5�����G�W� Z�{)æ(@b�����oo_e�&���m�=A^�j��,�5���J꧞[�6��x���יM݊dxn6g�b�]��.��R����߁�b'mI!������H���x�
�x�[��,��a���H\6d�X�����#o��36V�?��c�<������iE����7|i�ZU������/�hDZ�5�5��{!���*�~:9�
���g�G/���qЉf:q�K)*�1֨�s���k�ׇ�,m�k��AӃ��L�sL�� ������Y���(9uy/�@���$�xZ��o��~�t2p�������ŇSx\�Y�b�L�q������ݬ�_�q[-�ѐ��^eѡ�P�f�X�o���5=$q���DyJM�Dۤ0~�9�"	N�;]8�n��=�Y��=L��� ΅����ƘD�˘�i��k_���M��D*�~����T� �@�H���,�5��
M�L�0/�R�X{�ҕ�x��6�o �/�Z Ҿ�xױEw�ݜ�؍���#������0��-&�O��!^gd�ә/@����ew{�oI��V��M�p��d:ߕ�Z"��O(~?R��x�!�t�9��T�QS�*`!���@����L��$^�� �7=��et{ڮW�t�ƂO�g;%�F,�A<����)x�n�!5!J�(��S�*!��:|���^B�g�	M��p��zٛ�~Ҍ;�(��g	����ɠ�H��6��Rٻ�]d�8���Jm
��KR��u?�Q\4vc�q��3kxߕ�����L����_�o!|*lO�A7��k�a	���&��b�m�_���`W�e6�jv���4�V�&Eb-U �����'�C̄`�_���܎���z�6
��x^2}�r&���vE�Em�uA���>��KH�C��8"�k�҂�O(߉/@���DH�2� 4�O;y�#l���Țzŏ�o#[)5��Nkϓp�Q���	t�g�q:?{Q�����E9��h%���q)_K4��3/XK!�+���߅��%������^4mk.G��b{���AޕW��V��a�~�S��k5[�Ж[�w�����~e��j�X��R�o�^���7M�(295��w���4&�0���2b}/#z�4���F�X�
N:�wzL*����{�vt�G��.��xP�3j��?��ʧ�+� T#R�V�E�,�_���5�����_���UA�{[G�����#�J޳↍Ix���n���y.�%g��!s0���X�Ƙ�$�?�J�۠���D�nR��V���
��܊�1�y$�$W�Qk����Q���d�iaq���𹚲9yL�5�Y���}���&sd�a��������y�9�<�z|Fvpׅ�(��Je��!`�*�
�7��2S7��T��^��*���w ��&&��е5�H�e�>��Ђᚥa�O���P$��"�O�mV6��[��뵤�W[m.��	R��
EQ�ҟ|5� )���}�V�Q,���6>���ņ`�Gį?ԡo�i��%��x�j��el��df�B��6&ŏ)��c���9�๹w���;�KD�<ZD��+d���Pc%��e�}��w���Q N^��f!^_g��s��
yH~�kZ�	|��i>K�ɕqR��D�� ��4z��0���3	� ���
m��(��8��$p1]�A���+�H��7�$-!�!����k�k{����ɔ���.5(��l�'���{<ޅ�	tqt����'&��<�୽�Ar�ǎl��dJ�6X@�|4c)�|�(��C�d��,�����B+�O��ݔ���o��o����v}�Jf��7ڿ!Ú�-,�p=�Ʋ�s38�5(�g�z@�QR�F&L�0�I*�S ��ȥܧ�����=���iU�O�@JE"�>l��
���w��V	�6�f�Йގ�n��'��d���_� Z)�������YO��va4'��
�Da���qӨ�j
odA�_cd����������L�%OΜ��!�yV�.s��\KP�R���0�����z��6���\�g�2+��A��}�A`�v趾;�:�/�uC��E�Ϫ�%���Egg�,%^<�Y�Zp5��A=F9-1�粂�r���1�A>")L�kp�Q6-��DTʵ1�L"�lizGG߰nch�*H���u�� � 7�[��uv˥�*�9"�g�}�����=7$K}V��}>�[n�6�8@ƭUs?��Si#&�M᷌౅x+��z?�����,M�V�`���2������N`���}�/C([�p{����;��.(5��j���zg
M�������Q�iO�s��U�cN��%_\]ղ��y�Z������m�pGX,�T���+��\��푏K�������:����5��� �ɶ��~�Q|�Y<��ג\e�_W��k�w�e��Q#�O,�z���=t"cs�93�!��|���M~�m�>��*�U*	��N�L �Ƌ�k!��͂���x�LH뽫*`W�h�Q���Ė��Ue���+8�;+5F�uM�,[\<�s���@�8�(� 6�Z�v俔x��I�R�.3`Y�Gv��
y�-�&�?�~���d���2bK�e�8#��Y�_h�|�e�����X*�dml����p���GL��ucq'���[k�i�7��	����ٛA ��Zy8@�3����� �=��q!�
ⷤ5X��h��g����m��m@����	���]?��1̪bL�'+�Vu������z8z�iϻqŬB>�z��-L��pK��.S���~�[/�s}��_��T%/(Y$��u�K$2����:B�� uޕ=����!���EG��H�����./^#Z��
c���mȅ�S~�q�kI���Yzy8�o����s\O��y!�Q�ͤ��Lm@�K�\ş/Da�C �����֬(���AcΏĥs2�IJ�Gu�B{N�Zc��AM*����&g.m߁��w��S(,��^	:7�B�kaT�D�3�ʣ�䲈�F���Ag�lQ�0|B�<O����(��ё���8�7�ֺ�ާE.��s���1��,zp���~��ZB'�)��QT0��D0��p��2�q ���ĭ� �b"�)C*i�t�Z�t!�ףG�J/1i�qx}Rb���AL��r���fx4�i#~��_���2��SYF�N#�	1xe��(�e#u��>�o�0M�!�8�C�^�~0I�uw����7��Bk���-�;��F�Nr������#��fn3#��öK����Ls7�69���O�$Ղ���&V���Ἅ�`W��+�׊2��1?.9%���|S�;����G�-�vW��{�X� j��<%qLM�E�T�i����Q1"�0��]�����6N,��D�_��O�R�ս#��}�)�>4q'�5�-!�(�Y�_9�q�x��i ހS�&	Tۮ��gZe�PF)d�B�h~����K�&��+j�^%|�'����/�
4yV�΅��(�wX`�&ڎc���?'�[��$)��6�,w�̈k�
�5@��r���}�����N���Rv/��$�Lo:0Q5�"�N942���2&Rhq߆B�C���9��A�H�����Ok�Z�aЯ#/%h&�䮥dC�B`�}`M�x�F�h�et�p8���P��� ������G�Y����
,m����P ����S��i�/�b���x��:5{����R�k׵���'�<�w�`p��(J�-*;���9�݉'�����:�'S�X�9�(�s }�No�MPp?��1V��bp��W����6�ȍ<D�_Y\��ʔ���5���v��*UV\UҭZ�%��$W|��wUɍC��Y�#�K$m�T�ڪ�����}�?��CMr��7E�,tq�a��\	4?r/��V��vx�X7�vE5������3�_����y�؜�������H,��x0��=P�Hfh�g!\ƨ������Z��k��@����;K��M?�ޮ�
q�0�7�0��^�A+s�U4�6��vk��������s�#�J�6�kh;:�P�^�x%�Y�U������N%��LalA:��>�O�l��]�(�%���gX&T�1th�|II�nx;�ǀD��[��(�����ƶ��6rC���0qw�hSF��	’:�L��m��2{.����Lm}g΍[v	$����2�#�⻤{�mĶ������ Gѵik��P)'O���˽v@��Y�yT��-#Uu�u~�-4@z�)�b��p�m��q�`��KxH1�?^�!� �@\eЯ��X�Ռ3���FX�"/�����2�	X���܉v:���d��� %�"F�j?lƜݱ9 ���P'�p�� �SlR�sɛT��|3#�	e]<na-�<q��^Ͳ�%�*XB�l7��-��<�\������4J�_~3Q��،��N1��7\,��a���*8#���hu�l\�)(��,�3�x(iZ��iP-k>C���Z�A/{u�c_}NU����� �f��߹�'�e�b���T=&���ָ+s4� �Z��q����^Q&w��a��H��UWB�ϩ���-
f´�Q�}��c͢� גK�w�2�e�D��0%\�"1eY�&M�d�a�1��}@��e�%\�Ib�޿K瘵e�'=F&�uA"�ܗ= �����zֵ��N$;����Ծ��8 z�R�k�D�|�� ���̆nŮ�+L:�b���U��Q�����\���(�����[�_$p4eQEƐۂ~!2��z�:��>DY��to�V���
�=?jN���O�(�@����+��_�ʍ~�A�Tρ,����<�z$W�4�.�V�i���fF=^��/f԰��
�@��ՏIL�拀�2����$HR����Az=f5��[uJ��?~7({=� ���|�|�}�m&$H��G�"���P�[no���S5�9����Rfiq�