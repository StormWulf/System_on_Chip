XlxV64EB    55c4    13b0�Ҭ'k7�<�Ül_�W�5p�m:��W��fwF�U��hR+�T4�����ABW7��� {8�-1H$	.��H��F3�m��k�=��)5��{�&����\@�� �+��|J���g�V�ט3Á����ԇ5nJ�WI�ӎK��2�pt}�{!./?�^�r���v,x�L`)��_���Rlt�=C�,�G���;�`����o=d��^��E<��,�9�DۖRl�1MѠ��ۆo��+��vCI�SL�](EI��g�0�R���{v<��ٌ�%�F�`�'`�Ռ�̅�l��ۼ�|&إ��^ۯm�p>
#D;���.[Yy5�	=�o5�����ս�0��,���?&�:��޴a�T�t�k��=D�kМ.��RWvt-I���,w��Y`\�-��i(	�v5���#��2�âlڬW%5o�]0�(x��$u���5�ܭ�;I�}_6��,|;���It �xlT^.,d�|t&�_�]T��!#OP"�9�8)���$�:ؗm�����f��IR�}��ܾ�+$�����f����7ˇwT"O3�)2�����n� �o��Aec<#vN��r�bĔ7D�����t$8�?�1��w��_��]�����6+���ϙuw�^��g�B�Z�N���{H�%X�F�0�~:�9��Ծ)�Z؇��v�_��8תa�8'��d���A��l��|�W[��р�Pj�ݧ<�FU�d�`�ߴ���)�h �uL}��ef��A�j�+c��i4�+�y>�G ɻ�cmc|�S�pY��|�-��.i|,L����j�~_�n����;�kg�"s��k`v�C`DjE�s��L�|��g9B<�v|�����������n�w����z��|C�T�|����rmJ���X����,Z�0���^ך���Z�l�L��N49�%Q����r��|^r�*z�Ǌ�͈��ףa6����l{���s�9?xZ�L��5����
RHl��IF�����i��GK8��#�d���F��� �ËM:��;D�������Y6��{�l-n!Qk)Ɣ
|v4r��/��w.�k
ER�ft�KuỴ%*<�.O�b��N1[sv���C@�Q�aN���e:�岔/�<�fQ,!Zp��^�hT� Z�g��g�Jə6�̈���G�T~������!��1�9�0B(ͣ�)NtE,yM�ʒ"p� ˼4^,�X�h�8zb�R$��8
�7���fQ��H:wJn�Bٲv|�	H���c��@�=��vgԱ!�E�PY�AY�SHU�t3Ch��)�R�q�z���˾��Tvp�yǨ,��0Ֆ����%&�r�c�@��Sp�]sH�?5:ې�а�p'�����(�.6�!���ʧԿ� H�T�>���%�˥�L�\��fl�|�ۤ�A�7�Qċ��U�<әۘ+��.<֎2�.��'m﷙ud��k�ik\�P��}[!V�T���-w�U;��7�!����ʤ?Q�!�
����VYux`���u���Jw,�๒���:p�p�ȡ�~�ًM���e�Ǚ��"��ɍ���{1 @�/����5�(�<���nP��j�x�iNc�$��D�յba)�=��%R���O�/�WM�46��gX7h���'��PҍR��*}�߶#�����ʑމ�Ě��p��#�w�5���5j7Ӄ �&��%*��$俪��w����0­�J��.�tP����~LIH�����7)�O/��QL�GE֩S��.�fq�թ���
�즻k��y;^,6j�5ܯ�"��$���5�p�  M�e�D���$ꖛ3k
���+���13p!��m�d_L��w��T��g�Z�� ��ǝH����oqjE1��4߉AI@^n!�( p�	!�2�7y
��'��3E��Y������Y��p��m_�V�y�J5�AE�d�^��<;m���rM�3)����� 8��������籬�8��fc�	t���łōY^�������z��L��G�P�
�� ѡ)\�B�d&?IW�N\e���V���>�÷���������r������=(&�̿=ĉZ���+}��;Cf������>o�~0RIz��[��]�H�Ru�yO��*Ӵ���H�~°�b�x��H͇��`���c�� gU!�C;����s��J�?�]���6|�v�����K�4L���c���8v @-�#�H����Ӄ-Q��;���X�D���� �#�q��[W�}��P��W�T"��9jk�\ya#e�����(���Ͻ"ה��Op @Rl^��ނ��o�V|>ϕ����Z܂B���E�Il�EP�V����I�<=���0��J�}�������y�p�\��bE����Q��H9ߴ���Hg�������~ZQ��A�;�Z;3t�c��� �1�)|T�K*��q���W�^=� ݚf�+��~�$��M<�r�Y�
�1|�\-p-u�z���/���AV��E��~��B74~�Vg��e*�v��`@X,	U}yJ���3�Vz<��`܍:Cd��P�[Ƌ��r�j��do��t�,Tt������Lx��H�*԰��|Up��cCROf!^k/"���Uͪ:�C���p|�Q��h#���N�QS���Ʋ�54h��;Ni����%����TV���s�mD?B���
�1�ѧ���x�l�̹^��ipʥ�[�<³�+/�ĕ���--y���g� 6!Hp"�D�R�O`y�Q<$)2zR�x�B�}��'���p�F�0E�� �R���$��`W�鲼�$A�'�e:w�K��i���'�e�u���|�3� (���N=� ���d��$ �ݲ�D��m8:7[E2w��;D/�6�6����r�ao�ՌH�ɤ������7�F�-l;�����	����\�� D���K���ܘ���M�:Ǉ_�,�5��W,��V
���ҿD����g6-a ?c��E���[=o˘$8��A�g �l`����?h�L���:.��/���6��'�c6��J�#��8��o1�±���$�I��8���4��(?y��[��˟a�J=y��5?��'��1 �Ր.�)����K�<��oLTy�o5g�x����5��
�iYQ�������#:P�2Z=Kխ5�jf���=%[�����YU����};�i�i��%6��_�i�0$�9��U0S[��*��.�J���A�p3��R��)8D��7�(��^�"�S0�2���/��ߌ7�����q�{%���ʾ��H�ӪR&��a~7��Z.��Ż2��&@-��h�:�G�dA�LP?�ׅ�ZV���M���g*Ӊ�5��UJ��n�K��l!L��h� �χ��)q�R�Vw��Ս43}�h6�<L�o���3����?�7G�{7j�؀���n&�$X�ĺa=(�P�n?�Y�����y%:(u�f/Tn�}̇͒�>vS�����	�&�~Gj�7�0���0{Ixwn"�Gʚ��3�2��ŉ���S�"���]���a�
�Υ�`�AGb2J9���y�r�6�R�p�VSu��E�>=t�uL���,��!V!���4�/@�J��t����G�Ղ�S"<���ar`�ɜCc�%Y�������9�)�VȂq�)���0��d��#D�Ha��=�����ȕ���ݖ���� /���s[���������>"����Z�nMҽ�y��1v��U��h{�/��^;��a����Mq���D�To��h_U����<NK���]��}xc���*"B�1g�9�gѧ�l�A���}/�:�́�zJQ�m��#!�v���21]��/���Y�ԥ�{T�����/�6X���vv�:�'�9�J�b�2G��	,()���G���hb=oo���ɝy0�z���@�S�2N乀/�t���dQ����r2B�f��b2^R��	+�����o��ƐסHz�x��As_E�e~�LH�8b�n7/X�08�}s�����5�ǛqK�ZڡՔkN����-5kR�>�������s-��Y6"�l�Q��������5���Sh�٠?Q-/"�&��s���v����H�'j^�F�����NbӞCS�tZ&,?�O�����FZ7���**"e���w��b��I#���:��]j͉���=
�c�B�ĩ%4if�"#����G���_�ޯ����?͹dɞ	:|[��*�ف��-�w`� ��K$��ƛ����q��(B�e�'���47�P����B��A�`Ϛ��]U9¨���b�F�S�1�����do��� k5�z��\~�@�o�I!�8�1(�v��E��uF�y(��`q���b*і-g�w-2o�Vl��Q�l��:�ǗV�u���RE����	Ne1��O���P��儇���sJ�4�?S
r��ݲ����0��J����.]�������\$�{E w� �ݹ?�	�H��
~Y� ������^��ͨę4���(�������ה�㖘4�T�?�%p�=���Ʉ�^  :���m$Kd@<�1U��/a@�s���f�#�N��\F}�(W����;V�qmt��cx�p��k��H�_�����\:g�7s[@��{8�R�Em�Q�����oS��[�ͅ��X<��� 950�G+G�e��a
F<�9`̻͊�{{�>˛� ��M�v�!��I$��u�g��ིq2C��f �X�e]�D�}�)6�m�GF=��Kƨ۫ɮ�ݽ��A��R]��yV?5vĴ(��9 5�V�e߇����ZAV��	���nS���y�Fȭ��h��\��|ﰍ���$�WD�F������?�lҧ˹����}��Q�4��J����┫��4��mua�dumZ~#����燅���?�Z���b��{��<�f=����I�z%&����_+ �S	4��+m�