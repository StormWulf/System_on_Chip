XlxV64EB    589f    1210}q�_u�v�D���/:ɔ���B�Թ�0%w=����j��zIؐ�[[P�ۄi�d�;e�8�h��)r"KW0���T��'6萍\�kX"�}�p9���a��|���J��
G/�qd��|�>V�߅��֟|̈́l��u��J��P��K��yտ�̲���b��"|b�YKxJi]�đ�[)�rUK�e��#l&p�n�$Eu����O&[������V���CB0���k�w���)'���P�
IB�o���B�`��搖��X�g����B���aO�)�������> B4\FrF��u�@:��'n���x������<ށ�r��Q���Js�����hr���?����}r�4�<�#yy�\��~�X�f�ʐ�j.蝋PzHѬ�r�*)��+���֢��S՞Ր��y�j�i+�9������o�`�8�I|��tA#���w�y�j����9���l�F�[�98��Fn��͵�E�)$VY��]�������I� �GU1\B�RG_c�ʒĳ��w7\�L���z8v�o/UEd��l��, ȴ`���ce�)FM'5� �9Aw��xˎ��f�@���?'�����@Ϩ�s���ɠ�}��hNp/dv,o�L������t���J(��n;�$EB��uC����F�л�0>�(���D֓2+o��Jի�=ݖ��t̎��))_4|Ո4Cc�z��e���M���'�kJĕ�?�@ڷ���4��c����D��WG8�\�zt��.x�M�-��*+9G�����	�9�2\�����	��N/�T��nUN�˛���>����{}ph�i�eUǻ��aɗ���I��]�,4����y�����n	,��Pg$:GCP�I��i3��xW;�	�ꓻ �{ĳ
�7�K���B>

�1�O����w� c� �P�g��<Utw\)�g$����7h�֟�Vx�"hb���j2RD�Oْ	T���D�t,�bs7
u�a��v���Ӌ�U��C3�������C�Sɦ�no�u+�G��F�������c�0u/�{GW��W��P���	a8�t�2��'��Z2�<�;]�O:W&^�y����һ�X�뉊����T�Z�ЋmH��~��J徹��&�-#����/�]޾�nF�5u��{�� ��*m3�*���|�ofz@He���)���@i�V$���_��nD��|A�4tŷ-���6erI�j����x����H���4A����CU�G!�f�U�w�\��Y�p�q�4��V������
��GC�Yb�4S��U��L�q�`v���d���n�
��#B��A쟙C����Dʘ?�1�6���S���z���o|���3F�B�f*��K:P�|�x�Ǟ܈i��B�<�i���sz�6��]�5����K����T���L�jUiOQ�[�-j5�������d/��p�ʇ�$�T����WMH��#�F�����!;�lU�nTӸ+���w`̎�<���@2w���>��@��҇�>�t��YoE�{�kS��!�!�rH��HOlk���[���^�V�?��N
z�*�*7xn�E;;d3|Q�X���\{Hl���t5;c�vCT�?���3�wTM߮ Kl��~(D�ݙ���F��tF�Kp=z2lŜ `�Aj�Q�|����\{��}ѳ��������M�D/Z�:�ﳖ�&�S��:���SjƬ�'KF��pIe(
��I\ɘ���,\�7���\3I��gu���m�r`�7x��@�Y�e<cl�d����M��T�k����ŧ~�D��f�z�a�KݨJ����쟖�{av$��z�
�ذ����pOA<��fE�N$�z���Fˣ2��GZ�I}�����*��Z�ݷ�U���UQ�9��}M�Nrz��?N�|®!O�:�>�����3�䒘��Op��=��@#m�f����{�;���lڨ$�c�aԄ�86�>x@�9y�v����r���6���8�|	^�P&4�5��bN�t��=6�������*[F?���l�%`3�Da�A�=��%�`zrAa.g����D�~�	����C�;�m�^����Gr:@jH�|�,�լ$�_u(�)s�7���!��Q�Y���P|���O�܌�%����'n�G���0��e���. ���,������;jY�����d�m�������r�g�l=����\��>6�j��n�2�1����|@#��d�;z�Z=Ō���=����떰k�p������4��|X ��N�|b�� *�þ�yQ �\b._o�Y͛t��	�𰿚�efg���S�4";@6�m��O�T6���#�O�����Ĕ�Z�x�1�k׫���8ޠR�b1I����a�s��/.u��{[�["��'��R7Mz^�"�CAc�&���~���V1ǣ�XD��y|�\����L֩�a{�)�~������?�����Z-5�X�N��W��������4C���j����=*�A�RV]LXUZ�s�z3��ִ�� 5Y{^/G6ͩ��R�:J�Q�����
T���irKf�`�!rÍu���j�����%�z7�
�����xe�\Cm�� D{zy]�@ܪ����_d|'&��\,��!�1�4�$��;�Հ�ɵ��w\���+R`'� i�V�ȫ�E��I��hw��]��[%�E���%�_���=b*�.�YQ��#KY�z�<������d]j֩�Ł�J�#�4ߴS�MS\��X�cys�X����x���?:��[?�"�;�NP�-�n*^[�]�L�u� "D{(�A�Ce�����0KĔ ^3�F��Q΍�^�C���#���MJ����&��$�!���)�y�z�|�|�=}{�a\Y`�y�*M훟�L@��N"ܞ��_X�/�+�k�Ĝ�>M��T��<�� ;���Tz��q��%D�JN�����%�`@7X�fjIZǧ3 *����`�}��q:�u������E���AW2Y�)2�[�;ͅ��=�*�QCO�9j�x&�m%�k��k��2���s���)��0�}E�Ԅ��sW�Z��+d�~"��0
�)��d�Ц�U��OF��t���д�L&u����5[rb�nu� ��'���������mE(5���s��G�P��skg��0�Ҹ}�"w����g}aiܘ��Hc�<k�6j
�Il�o�1KHH�����Y58'2����L��]^�a�\-Lօy�_@B#v�Y�E���hq�H
\qߢ������o}mD�f�X�0w0Q!#EKŖ̝w��p�ry|SU���B�����Y,Ь�H�=� n���)%ܩ�6��Bc
��b{t;�e	�R��ߐ뫴>S�L2�ȻJs`��>^������"�e�%`�s{�.�࣋`B^�H�KuU���,N�,�.�V7��\8&��@���L�;W,�ԪL�0���������F��7LЂ�v���(�ת�g:�c�rF���.���_��O���v)͋k�]����+u���<d�VK�E��8���7��;d�Ora��"��{��Yf��ϼ��Hȣ�"8Y��̛M3�2���	r"��V�e�5�>�6L�����
1�fɄ��R�2x]3y�u�͆�
"��%I�$�+q�h��%f��3�'G���p v!n��i��T�zH�MsR��G8�i�<��9���	xu��.@K��8�F�U�X9�wa_0��i^Ο`Z�#5��w�e-�tYlP
%�~F����l�l��ȯ��}�_w�a��AM8׿Īw����EK9R����"�[�+�"9=ЯJ�U\�K	X��p�^>���=�O*�J���۵� ^H���� ��2k���w;R|c���:�A�fS����,�"���h��z����Ю�&��]Xj��CO�(�7��I+���̃ �#�y�i՜S�Z]Ew2��:=���.Cj���� z�r�:�d��H
<���Ͽ�$T?�F��.���v��7b�c\�;W�&̯ںƊ��������ʬ]���)�:+��41F{�x������-#���ڊ?�z@��T��;��v�1�]]���FR*}���i�2��"\�wգE#���"��:,�d��j�I)�u�iyR����(Ȇ��|u��**������))T���u롣;Z�ewUm���_['�j�і>j0AbXX����
y�Q�(�W�k����Q��h��,����FcY��pB�1������v����l���������7/���Or�)Q�j)�AW�W����~V�*�4��L2pͮ�^�n[��u�I!��)I���SĔ)⌆���4��P��'�+K�<&%�1O�Z]L�%h�X`]�;s}�e�0y�⊍�#�����f�t���YX]*�~��>]��\C�y 6�5Hb�~�M*��{.�T�5�!$�A�;��VB�}�1Viv�#B��k~a�?v�Y���j��h�2>@昄"˫ ���pr�I�