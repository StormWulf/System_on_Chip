XlxV64EB    31f9     dd0X	/���Hl0h=d<zw�#� ��N�g�0JpO�gh��֭�q�+nQg|���%�2��!O���0�I����#��6��ck���_|��"o��?I��<b�Q�E�W�6�#����!WjZ��9F�X6�'�ȯL��z�!`����Tz��y�l���H�?��@x���)/�1
Q�t����6ٔ���|�����Y5��b������o��39dX�9�7h!\��p/O۲�q�{��i��p��g4S�"�wLx1&L�H%)ڇ{�'/��!)�4���u�^��ߩD�̘�|@FU��:T�����Oǖ�V�3v|Yd��̕S=����3�_ H+.����Ґho��$-%��}HO��n��(�C1�JH���	��V6���Iyי!wH��P�Q]�[���o.]X�.�;g�hL���O�
���.��B��^�V�U���i�i���S�M�-U�c���`M�>��p/K�bT����3�� ��c�點��%Ʌ �K[6�4�B���-}g6xndĈ8vy&z�S��!��Y]��t��l!^=�&�VEg�q���<����h�$�o�
�3bBX��V��zu��p&���I�����MRY��� �pΟx�;"VtBX^�����D� \{�`ˏz+�,�.ǃU%&�M�N��3�<�����'�ju���Ϝ�������K�
��\����Eû��g,y�3��������R�G%��:��
I��R	�.��{W�r�#<�������dU��������G(��,�X'�)�ԩ�t_�"���3F��vy�)'�mO�v���O*��T�<���ys�
;�d�VL$Ư�vŧ�}�����,g�&�]���0�m�k��V�5*�ޅRGCf3�x�8�rӤ��L5݌|E���/iM�;o�C
�R�:�#�Y������2�\�]���./��X�M��C0v��n���=1􂁧��2���ɢy�cL�-T[�)䂺����B�x_���H��hϓ�(������(�G�ç�?��"�����`�(��ǎt����2 �f��^nrZ�H�p|�	?�`ҁw�1h,*� �fUO�`��S+zb�G�
�ڒ�%�]��h��+�gǵm./�)g�	��fKL(fz��������-��:5��+�8��m}ylD��cș4��]�5C��gvV<ƊtF�LrH�E�pSX�/Z�!�����O����'���V�0��iݐ��
�׀u[5��n��vt�a��tBq�����7�����}4/�֏8+g3/�H/���ɯ�_Od��_�Љ3�Hµf󈾞þi�9��V��>П��#�-V��:�՚*}�d���	(/|�L��D(t�4�2 -y�BDO����e��&d�fx����(��l��m��� "Kq�%#ߏ���J��>G��k��#���K���ʦ�<�y�;��7������<�p�nY����0���	���RzC�o���ۖ�H��L_���ӣ�
S�M�� �����]R<^��֐g.@�˻�H��.�#TA�y1�rhgXRer
zS<_�9�2B݀�9�4KX���Z��ܸ5��=`�ك�z��"X�i����s��ա�:!�����/b4P�fZ�"X����O��n*$�Ig��F�����]ũұ�Ś�=��8���*�D"��D!z+��kl5쭟'�.Q� �'4���MܯM��m�M�o���$
E�}ÿY쳏�4�8d��fH��l%#U�?ۊFX�a��!����=$�R��cp��Ӻ 0�	b��vp���`X� �;]���?�jC�^p^�,��ȏG�n"�5��,�4�`.Q�i�IR-� �{��N�5�;5~;��ϸ�G����h��T�QKՓ���g�̑/�@�� �0HN��h?�F2�q��R9�n�ixeC�9��˼�%lB�l�'}�Iq�"�����b5뭸��:��Z
��S� �����]�߽/��p���|���8�Z�l�4%����Bݹ��yY~�������������J�e7���S�� ��S����,ݤ�RҮ��U �C��v���-��7@؂�:~C�4�ɃB
_��~Ql;@NN���E�^c��Rk�Eh�	�]�J��d#J�^[��0��������]w�_��T���ړ�
������Ԗ*_��=�F�<�Zr�	[{_ƥ<��/�R<޹Y����ٍ�M~�һ����y!Aq��sm��}�ϫ�xHf�p�:ڴ�	�k�M3g#Z�X/;w��V�������G*��v��cT[��{	���z�0��)"�"�^�w\t���� .�w�"�4�9�:9=W��H�ڼT�[�һR��W_C^1
n
����p'�c�����C��`?���B5�W*�w�ٺ2;���?u�긖��&	+{` �y�ݪi�j��V]5�_?�LP��z4P�l�A����s�B�uοS9��*�f�7^�Dyj��?>�O�QL�R`�\����3\R�LI�n�o�g^a�/W��a���j?w���l_r�]�愧�;˦��OW�a�KXU,���x�S|�>����L'�	~�"���h��(),Y�E��Z�̈́�y]����2U�9�ն��Cpq�q�b��كAI  o��H#�nK7�oj%���c&WLw��0f���h~T�x���ƨ�0�ߵ.�?�M���8h�T�rT���H� �S�F�	�>�����qif�@ME�)B�

-C>X�}��h��$�g]�h����hDDkx�3�� �R��t�z6�YB3_�T��NA�Y喝Q/̽��	Q!����9��4{C�11�I�I�XAW�a�m�D�'ɝ�	��$���ZNP~CG�}����Z4Q$�h'
s��D={ p!�]���X�P��	�ԉ�۫�!�ǦF&�Nw���Y����Y��M��(ܼ��/��4���٫������o��1��A~�iq�¡��i3�<�?�GFg�9��M�A�֣Ҁ�3�>�5#qa�/ْ��,�h��P`]	
7�O����"3e��|�i���&��kM��zڞ��� �^�>N�w��Lk�ҝ���m�s}�,E	��,�C	�ο�"��i�fnS"M�U�%�7�*p>ME)�<S��!Rv�0̦E�����[ܥ�E���y�"�K��E�QS�Av��<���e��;P@�5�eI��IFJY�щ)Da����|ӎ�1h3��ÓY�J���(�yp�$:�p]c�D��\���kQ^Zb��8�"�PP�
��#�|�,�f~q���.6R��bO��鏥�8`�w�W��t/N��r�r�A��kW\:�r���L�l�剙��\Y�7��m܀�K�d���4H��/��J��4	W�q�6q�C��:�WϏ�٨-�asz�̝z���me��qmrcU$�UG��md�n�p���ƨ��k\y��>1"ӿj���G����`�