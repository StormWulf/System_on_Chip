XlxV64EB    1ad0     9e0��7a��a� �`/�eI��{bk�Y��qP�~>fІr�#e��,�HB3J�t-d>��&�xӖ�������[Ϣ�~t�u5C�/�֯��.��s���ڛf��]��?���F����Jk��sz��#�V}t-U��=_3~�X~�v��z߳d�Ë,B#������I�8��+V�T.9D��VZ�w������>+o�2Ԛ@:��Y����,���g҅*������ء�1�ZC�F��4�b	��5�6<� �蟓�������FA�V��
CG�[,L��C��C�M�b{臉��:.͏�,r�^���@q����oY����?�ώ��	�@�n���G�h.��A���,�U��aJo�s;袦D��{��Z�緍3o~vl�[Yu'��Tپ�zs�bz�*C(���S/q�f��ױ���v���@�#"��Q+�t�3��'m�=��FX������R� ������0�!�q��oΘe���V�m�n�S�����<�[��I�y�=9�0��k��D�1|��bl؆/��8��w�.��
 PK���xM�J�PV�һ6 I��˸�',ڙ����C�1Ie�~jl�v5_F��n��y�.� ��xx�M,���j���&�Tӛ�GW�U�2|h�7j�bK���ʮ�H���׵� OL�Ӕ���S��3d�*k(A�[٬E���&;>���Q���=\'�7�_.E-��'W����C�|� I�k�*��%�x���xa�q�G��ò����y�C
u�8p���hsS���O��&Y���_����u��[V��o���#5�x����۱M�����&�"�+��=Dn�9
��aǤ@�bf5�h��!�=k�Q�=�Bۊ�Z�����k&�h�Q�7��L�u8��P%�>��I�["-�zi�)�;H����z)�L ��%���|U{2V�gZQs�c7At��j� �}̎%�YW���!��%�u��]��Ctu��� |�����?�s&�I�۪I�@U�����*������ZS	�H�s	\d�_������u'�Cz e��D�`�Sa�����)���6,JG��	N�&����c�&D �X�P�W�m/[��{��;��O�L=�2�'
��q��AO�=��G 8q��#9�	�ܸ;W{{��C����!m�8��2��nA���-�,�(ź�e��3��P3��m�Ft�'P		XESZ�S��&z�Ӟ�b�F{��[�R�����(G����pܝ�B;�k0�F���:������ �s�R���C5*0��%��K��:~�|�f��vbQ'7y�B� ����֤�.���#�%��.�T���S���3h�{{һIQ/���8%�|Y�;��E����_���p�[��B�����kp�oV�#�bU��z�E�	�e���"~��Y��rĆ�Vf�6��y� Up�����q����2.M��[��`\0��)qѧ���"�Q��t��D��t�c��h��v.�K�i���c�f��Q��}��9����Ҁ.��Z�8���ax=l����+�t�m]�M����s���������q}��lz �X�#k����ӢM 	�ܢ�lXG����w,�@�6Q;���խj��Y�qk;�h�t^;��8�)?�n����S,�,�b�rO���t�U��I�MTdO���H�rG���E�>��YC�P��kH2��d�:�!�Q��[�6���s���XX����--��Wo�䒨P �?�r/��Z|1��wB��\wLE�LH�0����oU@�]Q�\MQ��|y�C���-�ܬ����@�m�������P� h:���Ū�I��(����WO�Z��)�rT�x&���b�j�k&� ��џ���}p���4�#�j|��u���Nܟ]���E�{6	iС���w������+ZAh�����k���%Z�ew���#h����⥷4���p���(*������،kI�Vb���<���Ѹs^��8YM��s���lg�}o��-��'��&��Aܪ��X๢=hޗnFѽ9<�ɳG@���ȅ́�äkŲШ7��j��a�6 �q�,�2y��ъ�C}PK�S��QI/��'�ߖ�G5G�f)y�Y��U��5.��D�z��6!�@��5p��T��bSp-���0�q�A��m��65Z�-����|f��9
�]�lCp���>+��ŧ_���Ѿ��I� �-E^��h�`�-o�tf� �J��8Y.X��Sv'�En�l�/�^��O������?�4E�>5��i�&ʊn߭�ח
`9�*��������k�}lA!�L���ҭh��\9�}�g�Z���x��PHI���v]Kf�]P���t张�I��R�l9n��_w22��Q�o��EX��@A]r'������$��t�+�w�(���T���~��{_
�r��]K����