XlxV64EB    2121     ac0�� JS��࿫k<��o�Vq�c���,>s|����ZpG��s*6J��x�����*}!��Sz}+y!*�0aa��Z#/L!0XKĪ��@f���7�� ���J�X�����ş����k\9�ɻ���T2�%���kR�����l�;#��V���P�t,}�N��������m{��v,}GK����ÝXC�-��xg���EM����Q]�D��}�DG�d�5�� ����v��S��u�Ǿ�-�x��Bg �c� ��n1=~��,@)��'�[h&���|ݠǌ&QM)���
�z]82~��U��o'f�>ӻ_����R�F�U-��0l�A�S�v�!�2FۇI���>U_:�9L��.�=-� ����y�_�IӇX�Y� N�Y��~DՙR\V��w�$��?�!���(���85��"*#x�������VCc��qB3�!���3�E�?9���TPz�[Z�#���@�b����� ���rp�-X8KJ|7Q��.z�۾�:�F�����KU2Pp��R1��/Zxs(�϶��^�H����s�R�wWv\xQ|;v=b%������E>}� �7�eMm�IȞ�Afa�a�װM5q���n5:x~�O�:j�p|{̒�t;�j�?�u��R.���l�ݶ�xal�>@Z�Eg ��C�EZ�(��ӈt(�
[slڸ���~�o����3�@���}��P�/�� �$�?ב��`j�{�$�c<��[���+4���NF����}��pC�7j;�)�ջ������U��S�u�>�c���	26ޅ�N'd�����ڝeCW�\7I�%\�@��_����^����<�yo9V����<D�N�ݑn�c�D?�}<�g����LVNU�:�xP�PY�g^��C� � �����K�]H}��gH'�q",0q��%pD�AXWo�`o��O|���Xm�;�cpD��<%F��ζ$��E ��?�6�8��Wn'Lk���6KB��\��l�OsB�L���6L4~���D�o�@�Y�\���fZ�6��kA.�q;M��M!sP�u[U���#�SP���'�����}x��2��A/����ü�dX��\/���\�C�	ǔtZGp�Kc���3�2���w���{����dek؃J*F�HW�~b�v��r���K��x�%�-l&,ᯐ����既M#5���ԄU#����u����p��[/����-��v��؉�tF4C������f滥Xf�]䫌�GoTv��|u�� �d3CY���i+�����W#�rG���`M�0��I�(2.D�fK��5LJ�%z�ۃ2��*(Z�<<y4��`�R���}�Mm�ㅟ6��'�Q/��42��yJ����)�n9$b���s[��.�!��n�O�oƹ���:��P�K�� �՟�x9�Q�?{�������!(��a�	�Q�Z�U��
�� ��$��}^C�r�}ѡ�Wm��KG��w+D��ʥ��2��Cq
�����<\빉X�G���;�o�yҘeP�_{â�F�mVڶ��f�,8�b�����T����c��H��;)�6B���������e��^ͽQ�R���݋�	,1yP���*W�~X��g���b�k��̾�EN�vg��������VA����/����}���t��l��Þ�P��q�/���Mn���w�}*;\��:4q�c ?��<n��_��� ��ǄaI���0�9%?���Ȃ(N_j�	�A�5�3�5.��N���h�%n�9��y3i��?�6����)��؛�%מ��դ�?:���J�3y�}�雃��|��/b]�GS�C�����H�������~�
5cUvq�t+%�xy=���C1_��%��bk|��d��Ғ��LT3i���z̬ѭ?K��Z�{�Mp�}��ߑ��s�QW���L���4<�˄�uI��ab���YZ���|�b0��0�I��v\��(c�%4��q�Hϊ��[ sGmM�9g�e�@,�t�����L����ͻ
�~]J#�� ��z�rK6�$���� �0�Y��B�!D?3󮙠 �'��q��4����׻�`�"�|PcϸM�F���F�D��9lm5�L��aw�tM�G��k'���j�t�YO��!\�Dn��MtM[��sn[n��j3u����)%k<��%>��4w��vӾ��G�����{-Ȧ�@ӡ	�t�Du{NvMo�}��ocs1��2��m������2�d4dνx�����m�U�I�N��8������K�&��i@�S�9�+w����2D��7Ke�(<|s������h	�߳�&��|gHX�(f��%?-?.�?q;� ����������S�����o�e{f�u$"Do��/?�K���TWW�93z4�� ܄�S��y��Pe�h��{%����b?'�!%Xt������X�����o��p?%�D�ӯ��Xt���|x�� a�W*�m|M����}8o�GG�b�+����'��g�~<C�!u�c����H*><�8�_��h-��A��q���Ǐ#p=���8n�C��Y� �Q���E��0���9�3K�+7O;�������^�����2�oy]y[�D��h<^����g��ߍ��@ko�g[ z��r4CS	���]=q���3�9�U0���Ϩ���79�Q�A�6:]�n���!H���U��=[X�