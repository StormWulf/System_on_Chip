XlxV64EB    6ee8    16a0=&a�ycVM��|�,���X���Dy<p�(�����95=Կ;ȎZS_���$ᝳh��ܰ�����������ԣG��ٺؼ�sc��PM5E٧�`��|�۴�u��{������4�"C�+y��ր$���l�$K5,���W-��k�Ô��~���ٽ� y�9�l�'H�ė�o��}���XY���䭀�f�C�lw����`ltɇ�C?�>v�_�8�w���Y�5�Q5$�M�`����l#��+0O��<�E��Z<��&�%(��O��)�*�xd�8�h2'����N�e�ҕa@��(P�}������{~ub 8�V6����$<�UR���^��F�Rd�b�����>����eJE���gS�x:��'���s'䶇q^ G�Zf��-#C���d�#�>_N�
���7ab����/D�Wg��O��O���#ҩu�ZZ6!��B�x+ȴu�5n.����!��@G)	��|N8��AJɾ�E(N�/iK�<	+m�j}�5��sAR@|�d��,�;jE]�Kn�ʏ�sPa�u�>���ƨ(b0�,��> ��
A)3�k�\<��0�E�񵇵���B2�v�:��$�2��*�l�q{��1�m�Ne�� ���D ��!�hpL���@ȥ+�P,q���f��*����a�K@A����K[@��7������`4r=p2Fֵ�'z� 
�;��4���~�?s�'�T������Ŀ?�-�ld_״]�g�r��;���Z�EX̨�Fvk�y_{������'������T�SX�Q{�����\ұ�9R���]?���P��:e���ZY�7�:��ػ�V�O2;�K�ˣ���[�J�Ʃ_�u�ŃZ��9گW���h�Al��}+�e���Ç�E�"�&���5-bP%�����ub1I��Q`�&�r_%����TG׫v����zB^´����]��?�E�+7�hcg� �Q6dy	5h�&Pl����?�B;��AO�.0m�ԉ	9��!���r��
��*1�B��92H'��iźs�\x�G������㲑�!�����~��+א�¬�P���([�
޼�p�5���ѻE@2+%�i##��W�FIVB����C�̴���z.ٔz�>�~3p�&�M��b.g����ώ�^Z���Kq�E�\0���
w�*�%���P��Tj,�k#��t��B�� ��"Ee�.r�pE]PB��,-(gܹ��:3K�u�O����'r7��bΌGB
��<�:*�E�%���߇~���#S26%B�4�a�9���-$ٗH�	�q��τ]4�"���*����� �ց��� ��Ķ!,���<E�P�0�����pX- ��%�+i�U�����0s�L &��N�܆���e��|Q� w���ƌ5#����aILKsUO�W/����L��\c#:}U4��k�i����ߑ��pj��S����������5� �Ξr���͗6���׸�v���=@��1��e��T�}7dD�ܽ�t��s���ᩋ��F�Q�.ܑ�1
���)n���{�.o�I�/��j_h8��U��Ӝ�b=��[ԡ���b��I@��]Ь��z�]�!�Y@i�/���]� a{�LG�P�V�X��˷ů$�k[�at$
G��u���_��Bdw��Y)d_�N����-�Q�=��u��
�����W���ut_l�[��%�
���\W�)��У�O+a�`{��j����N�U㮸s�g�oJ����穧�\]ɓ��V؅䍁MH�?0�u�J��Ǻ����(<�H������"�n� ��h+3���=#����\��d>HY��AH��,�Ut��|P�l/� ,de�D�-�b�e%��:(h99�ZpY��Cg�!-�vN��L.}�e����@�$��?�j� �6���@�;�|߬]�?#��|�Y��f���L�%���!��җ��f=��x]�  ؝Ci0�v��X~����m���@oy����S�v��K ������S`�{(Y1d�l���x��lǐqa��	��7�O �e��s�hcb/��xT���z�y"�#�M��@o�E�_Y��s�i`>�� �����r�mVR�+������ )ܵ�SQ�^��4��>��$�z-{r��~+����kP��a�r���s��:������5�0j P}�B�@��Q\�&N�FS��z��9J��=`I΍,�i�{/W�l���1�1�Le(�	��.UsOg����%p�S�\	����qH��:lD%�M0�"�3k�^�傅J}/l�2',l�{��YE���ȩ��s)G3|=@�~���z�=��G!��`��Z�������7�8�0���[�[����γyVy����~�nT�Q8�֍����~Ȳ
� �
{0�'jd_:�uTU���L&�|Ck <�}ZxD3LI|5��9�Hs��ʦ���]��� j2\s�I�w�$V?s�'��~�p���̰YMm�C�G8n���S$b"��Իc���X����!��M�=��n�zY�Ў����n�S�-�i�l#�� 
~DGZ�އ�<��ή΂�$d+W�����P#]h��C��(�z�W�Kgٛq���AF@�8�E)�9�-�5����(��<�^u$��4�
At�2K�uM��!`<���~�S1�:��a���	�{��s
a��=}/�^���d��[��W�H�9*�2�ɟWs���i5A��\,���:�9��pk�0�\T���&\�4��/�HC��M*���!<���/��v�j������%��Ҫ�ke̗��:�S�<(:詑�ҹ��H�1�^�Ö/��+su�f�u��30Q�w�kHC�3܉�ܷ����U��'.1k�K|z��ͬx�n��T?��Q]"�u�gF� 9��tCj�|?a����3�(47ս6W�} A)V���	aY�V�ͬ��W�CA���Aԧ,^��ʕ5�9����:�s�b���1z x�����R�������a�e�xQ�[Q,)�����+x�,��lϻ�JZ:4n�
*
��	Fm�^?�Pä��$|dF;Қ@9���d.�����(�_�5�П�sxq�5x�ǝ5�
ΔÍ���<L���3���JE�/<��|�j%����t��ds����D��4m���6��j�I6{��d{gWq,ս�S�a"V�Q�9�-lo�O�T�{W��Zc�2�ɕY�K��Gc%���%����F���z�׍�����މ�`*d����W�>!�C���?��6���V\�6xΕ,*��Y!/��hRc�-���O�-d�Wv��+�J�3,GWt����a�nշ���?�{,��������r�<���,�`�r�fW����{9�ٞ`�t���]��ƞ�y��;�%%["�y�(H����G�ػM���iYyV91�W�o�y���*-�w�%3y�I�^F��s���XE�`|��j�B[.�0l���p�����I���p��;��@#��7)��;���Lu˱YI-Zj��#h ��,��ÇOa���l{K�%�_�X^��@��k͘�P�.p������^��l4�q��,Βqĝq_��Z8��0�)��8�X�@�ap&����G������V����+�>��b�x�H?p�Novد�䒼EU	T1uA�-�㌴����6�k�:q�t����\��u���e=�c��ܔ9/�e�>��5mY�K�Ě)��i����nB�J���X�mb�d�[qAQ
���~�S^l�
!Ծ$�[�g��	�<��Xk؍��̌��<:m��w�h��uڤ����mj;9��%�$�Ҡ�bXWW�pB1��n�~a%�KGw.��3���$QgN���X��"����&�;Һ$��2�4r��wY2rR�`+:I�d,xSYM�ء5��$�̽lд}3!Z�۞���o|����t��-��;0E(�_Ur�Y�f"�W�Y�����hl^��|�偫X��Y�ϢR�;�[Y��j9.9�ra<�A�Lo�
�O���VmY.��ǥ}N�pYT��^���
�C�M��ܔ���5�?czU�(�ϣ��ע��:	��m�!�!����>z��򺱘�I�I��l�Z(��nՃ-A�����*}O
�Ҕ�
�[�(� 	����r�����H~����k���PT ܣ%`��Un����`{K��I@k��oGc�@��U��q�f��ho�@���?Q�����	�P��J����"b;˭_J�tJ:��o�.0#@@�gW$	��L;�������c��I�T@�:�����E�ߖ�2�� Zd�V�f�� ��8��rtL,
�L�z�EZ�A�5d9�Q�E�}�U�H���Ng�w�fN���0���7�\�V?�D�8{c�.���qxc�^��͋oRs�>y���&����5t�'i�4�.�*��&!���_��O�H�Yl^�d�w�I0/+�5 -��#���~f�]mw�f0��f9��|c�\���'�|I���UO䧸HĲ�cL�s�zU�ӷ�(�,+�������-�;�ޡ�=i�9\��w��:�D�^0��t���~����kC�ɿ~���[#֨tR�����Ua�bR�Cw��L�k�P����%�͐�mm�Q�=T�����]/�^6{���b��.�PY�K�ʫ�0G�!Ȏ��F}�b޳�ӋZ���d]4$wz6߸�N>W�(ՙ}i]�v��o>�_[~����rD�1X`W|;�����W����A6hk>#�l��]��=���F0D��>�0�Vl�A�"���(�Ӻ�ڨ{��:��=��>i$^v�#��ݘd�g4H��p�E���(E�A��%L=�����N��&�D��z�k�dZ0���&��%���7�h3���H�ӟ��X�)]��C�������IY�S��S��:��������:��Vl�C�G�$O�%��UjE�-�B_��o�EC7�Ե���9��;�i͌�a�;��O��5�3�N�Sc�'u>��,��QI��4a,��A�6l�Ȧ�_j����,�+Ƞd���rr+|�/�;�U��>L�Qt�7�d"!Y����/��k���V��~��~�˰��io�^(b�Ζ��$_��a�֡5��#���'�+�#�SfsKOc�D�U�<��b�Ί���ʀ��*�:+����lG�z�p��L���d�6�,�	dX�'�	[$YiKݶ(���_�؄���7��/���԰V��䈴���9]�/f�@�oV{h���<�a��63v�s>��D�ڧ��I��Q:G>`4���%��#�V奄 ���R�&{F��ǢҶ0����Y	�p�2����h��=� 9��Vݭ�� *�H��k��.�����X<���n&�. ��H3$ƹ��������T���n���߸��jo�U-Q-!��7?��!�PeV=�0�l����5c�o�{2�q�"B:Xx-$��m��.�a�0Џ!�~�ЏU(���|Ck_��/ #��Ͼ��.g�S���P$^��L����V�eLݕ<��V��H�;�s�z���
4N>,Zf��י��NuE������ȏ��7�|Kg8��_E��O�<��i:6я���v����d<�4�Zc��#������$��[��w��'��0