XlxV64EB    c9ce    1a40�o���c	���g�,5��P �d������h
�"j��t8�:e�%cF�vJ��ʭ��2����T
4g�o�_ߠV�u�2j&K%
R��q�լ�5����&<��I��a�u����>��Ś=�*<��|yԁx��D܏B��>M(�$�ɵ�T��d">-}��h/��
��H��4<��;L�ܺ�m�l���uZ���6�P��{��F-���z��jX�e>��v]F�k�#��x����P����M7W�U6�H kL;��k������� ���ز�5�9��W�M1������n��.����yi�`�$�Q���O�Rم�/�?�xs��J�x�^ɴ��"����U�%Ft���q��䤶r����?#��*v'����i�ǉ����ܣ!f��~����'���ĉO��N������
g>Z��y�|K��J�_n6O�u�u�?�[�� �$	�%?�bR�5��]+�����ax��.B���3A�#�.�0�D�C��3��{�vQ�V�� �)�
����n�?��djx����4`9�Gd�>N�pԉo��Gr�~"��3\Xd���F᭼$HF�R"����p�e%�Yր�Iܫ�f��|K;B,$�
e߽�"�O\�����!V�G�'�8	�b�s�B��v�S���%W�V�Xvfi���RB�P�j��������mF�^�L:�\m���-}/EGXH;ri��M9��,��ƪ�I���TR���8?��
��b��i-�~���o�[��e{����PkD7�Қ�w̵���۝�L����H,O�!l?``���~uKH�4/++� �B����7��=�(~ $�����?�����;�hy�H��o|�㑮���wH��l��/�^�<g����;�&�xMM����`Zܡ�#��Ցn��@�2��!*��M^�ә���uV�P����Ԯe�~a�?�h9�r1ʦ
ܖ����w��;��mMet��9k�ӪJq	j����c�e��&Ԉ��1�|�"�%9=�d�>N,��p�:���!�Q���ºz���='�A�����ߡ���
�d]+	NU��Xp�bS�6�OJU �
�iź�/b^	�w�
.aZ�@r6�7��X�V~sFp41�q&K��W�� O撑���HO�2�p��^i
�P�U���N���SL���`z)�p�U�^�+�Eǹo�����*�د�Oֳ̬8*�G޿X���7:��5��"ҍ���-�e�_�9�?�%FX\�ZSK6eYܶ#��Rv7Ͼ5U?�������a��f����G�\�b�	��ɓ�t��Fky�m5��
��b�׀�^E^y\a�,�5/d��Bh��s礠��;�\V{�1���G+����P�
~@�f�=����p�T��ڲ�f��=�0Kv��@z��mN��|�{<�*ᤉ!�/"�3�f1	,T�Nz 7>�dI��I�o-H��)ݢ�q��z�'��(�/��+5=V�3�5�S���,�XЗC>PTz/�3��v豧`�&���W}'�\V{�h�m�}Ɵ����J�q���{Mz}�]���9-����]o��hJS�\i�Ci��WjA�M~���-�8]��O�OzJ(�G�6ۭ㗓P��6k��^�c�A��V>��ʣ�r#U.q��Qޱ��I&���3!��*�5.���t�=��UW3��~p+2��aS+d%�om�V�<���Xy>'+�Uw�y�b�VJ!t�h��;���4M�8"��i���Լ�Obe?S���6.4��O�W�6r#
��-e(Y-��9���&k���h���.>,�h"����'!]�?���	�7�<�`B*=���I�!�x������4� !4#"��"�ͩ��� ��mo�9�&��II��2�JqŲ�=&�{��/���Jq*&ƒW����{�W�t�"}>'�ŗ)�s@�ɵ�
V�V�٣-�����I�]?$��[
��'�z�M?pO���ݝ��j����l���$�L5(�}V�ڱ��!���5����b87岸9"��y�~��H�?}��c�G/����AM����lg���ǥ�Ǟ[;�� 1lxt1��y�al=,�,�W�쑘�.��N���[:1��H�M�Z���{�O�/��u�d"���,�8��)*�ݸ��9�z5�ƹ�aK0��7��B@d��=��4�	�$�r�ʕ�^kV��2�g�uq��������?7(��%�N���du����8��5�����AJP�o1���(ۤo4���k�`���W�j�K�"�RQ���'z�(X�y,vR��t0I<;��Ϻ�D�l�]ف��e�P�`��1'�+D��3�a|���2�`��z#�x�ԩ�8�p*"�r���5�c:D��@��\�n,BYD�tioG�^q�]*�y�^�3����8�j�f$������Ց���?qOq���#�������3�ȷڂ7�c=@zH��ZY/* 召*��N�:i����f������d#�1�&��?޾�l�}���mlC����t�[9���1 �hXBMRh��`��`�e0'��t�Q�����ZS_�G�"`ˬk����Hv,;6B��,͛���s`�ơ���xTj�9�ּ�hu���j.�������B��H���`*Z��d{����c1�&�N1C�ȯ�%[$�+@>��
�-ṅ7��V>	x��-�!��3L�׋�﷌9э�"��%��Cx�H�ς�-9��Wo�O����^��W�����2UZښ�>��;J{r��q��o~ׇ��pqw ��k�I�n�'��]�ܼIi���vzD0�_t0����ߟ%�C�N�Q�,����a���'ggלS�Y�Ѯ!v���o=�\@��E��Q�Fi���{��a
�8ې����	F9� G�0�d�jJ^��ʿM�������A�=#`�F�y�L�O�tX��6����n�%�(�Z���"�r0X~r��E�O�?�3�=3/��C	��5�m������{�m �Wy��?��^�'��<�x�s��n8�������[��Cq�vF�Ԋ�Fp3u	����dD�dR���E���%3�z���9�P����ڰ�˥׬s.�#	�� @���.���Cr�c~�%2�����]IMb���1�>_��w:I0ŵ?��%��ֻ~�<h˩��J*/��0�B�n_V@��g���!�lQ�T���ӶJ�M��95��7��Ϧ�{��McNN8�bO,���R�T��&=j&D���YȒ�L/_��>+hI3f�G�Kc�"��)��zdW3,輷��G�nV}��Jk��&����� M�B`�A�Ƅ`y)�D���NL$����RހD�jMj�run&ƻ�� zoy<V���b�K1[�w� �w?���9*�y�+s%�<����Gf��`��#r2.��_�t>VA��T馵�������.sd���ob��X�H�c���λD-$eRC�� +���[��e�%����m�n �������RS���pة�k�\lx��~�[O7]�)�
+�e�-6��X��l�N�ʲ����i�I���N^�5���a�U��.�mv7<��Oe��A͠��7�2l"���y����M(#6}�/�fR�G�N���ۮ��c��A1o���@P�?����)��o��f�`F���YRCj{a�3�gl�hr�rn�����-������Q�+"����\т���S� �4<9 w1�mErV.pR�6���Djگ�%Vuy�����!JE� ��:��H���B�;]h�(�%�:ε���Y���I�o���T��Xn|r�Y����UL��|�eCa4"1������*r��[��Q+��n[�8��hf�BK�|���O��3�89��_�h䟊������}���v�}8�7�������"�D3П���>�l
Z�]�_�|Xj��Z�, �eiG�O����[�Leq���tvpk��L�3���$yD���a(tl���h���z �0��VHl���1�X4|��S�;��9:���8�{�Sfci|�%h��u�)O��	���{��P	&ww�[�v�EM;-��I���N�n��9����T���#����0Ax*�^d�Db�[��)�e��("-s�띺��~�3I�5�7��XA1�|��z�d\n�3�f�����'�R�2O�J
Sa�|�ok{Ϯ'��z��9�����,��i6 d��K���MFk4���z����u|�c�Z\����������z��� Q��|w{XF��_~d���"|���m�Q����5���\U����"K��op!�s=h�΍	SZ�I��I�!&���RO����\���=��lP�QC��XѢ�XL�3��<��SbP���@|���x��ELMr��-?��<*]�{�7n�|�,�e������g{�䣥�����^W96S}7i�A_�;�����O���ԡ� �~JxFƺ�u�xT��	V��.{�z����Y��lk���?�X�g-����L�Mѡ��">��hw��0s�v����T��:#�)��q�%{��>s�g."k��pf�E`Gzu�#Y�/w�b�)�Z��o0k�M�������[b�UFÁ�_�0�=Q��V@�i�����xy�Q��y��m���0i��5�2G��[we�E$2��A�0"��4OD�Ƣ��sUx��A��ݴ�\Ꮝ����Id�jX�I���7?׹_����	�t.a� sɬ��׹1z�}�t@W����4����XYۣ�*H���n�ד��y���Ҳ��ˊ�~����Ujmى	R<Ѐs�m<�}�Ywq�������	��B&���4���55��@+�Pa@셧.1����rD�F��B��x�M��Q�����J�o�h��
p����yB��|%1�˝w�H��I5� ۰��tҙ�q�(Y���ї�Y�>������a�2�>W��KR�-�b��/.��>�*�c�	�/(�R�� i�\����\���gD���<:�B��O��`.g�9�T�����U�͠�FdQ�C�f!��'�u�^fmg��>{���??��i�c��k|�Y��k5��;��~�Alj�t�S���!��\��5=@9.%E���4q=�\��)��8+��}̀�y7�p��,�{�J0
d�̦D�|��rV@Bܭ�h���'X�|�����ɴ�/�"�}�@�]��=gDmzX��ZM���`�ߺ'��ߙ�Wj��9B�o�'u��Zc,�f�9�i����C��.<RQ>w4���ͧ�y�W��U{XU��_�0�U�y�3���H.�6���& ��ڈ_o�,\м���?�x�a%�"�s� Sb�>��p�(��n�Fʑ�w6/_]���ՠ���/��Q,^�N�X���T��k��_��]��íDpZ7�ݐ}�A�q��?.�Kͬx�����`�U�֘�n+�%��=�����*�
NUƎJ:� �2'rY�Cv��X��}�!
>
ч͚,��	,r�J�T)k�u_��y꼙xFZ�Z"Ťؚ�(�"'�t|�B��Q�پ��ہ�˗	���^X��DDx�0S䦽<uڐü��
�=��x�q8�S�W��֋���������-A�t��lF���&c��:~�g+�yu�-����oxNSd���1��W��\�j��r�d#�m��˦紇���Jkk��}~(|�@�w1�~p������WE�D��@�*y�$Ks�G�2<��jL��}x�$R�4��o��C-v��}�z?����3
9��c�ک�̝�K(А��^=�G�*<����6��G�=�	�a���}{��'/�y��tZ�M�c���q�ZV t�χ#d �C��sj��_ߟ/!Fr�N�}�d��Xt`2���vv]��L��H�Ҋ	3�8,/5����\|\ۯT0�{�8���*L�����7�QZ�Y{�x`���ܳ�/~�������V6UgRN�49xvI x	��G�-���:�K��������F��]m�#׹&��%��l7�r(S)f=�S�S8X-�˯ �L�f��c��K���}�rA˞����iFv}�a�[]�hˢ���l�6$s��F��8d���)RwO����a�f��EF.3�}���$^z��i"��2x~����I?x���i+�;�P���u-�&)d��f���l����)�0�eW��p\ʭ��E��H���Ѱ����)�'-��GoI��ZP�x��!�J�쌉��[
x������j��9?�Uf���'��>�����z�/���!3��-oX��)�3ή�S�Kp��1�T�����g���O�I-4ah�KA�Ν��͕���/.D
�?"�8Ș'���֏��aQ����PL�����uB@���{&Ê��3�u�J�0���V�W�,���@�r�������S���IOi�T�x���	�Fv��69у�o�㪤�OVr2M��]�Q����|�|M��u'Q�:}&��[@m� ���!Qp�ç���y(�����
g��-����@�ꤼ\*���Zݢw�le���`Z�j�Ik��୐C�Z`sxj�