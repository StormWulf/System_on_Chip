XlxV64EB    25d9     aa0B���9]�{7�h���d�9ȱ�|b��g?䶖	<:.��Do�z9!��k�b'a��O��2����`K�\()�<��f`��R{�V�㚻��?	�04_�YS�SO~c7��r,YC�Pr\V�m߶:@��:�S�ǏHˮ�W���3[�# za�U��b��>��9�uZ�f8�P|������&�-ә��8��ۢe�u�,��n��/>^?~�u�u��2�����rOjkJ�x�GEe���5�M��� P������ �ۈO:oT��̬M�N�s?h�jk�iZ.���N���;�s�e��|'�����R�>"$���y<i�pj��/�#i�����|�/T?Bi��4RS�^ڸW�ׄv_H��p�Lꛭ\ )��8·��wx�/O��6���kPwu���|�v�lT�)��i��X�Z���:�����V�t�ڏ��^��������m��/���x��O���E���	.���e���MiL�fCkrKcX�Q*�[6���گ[� }��!ޔM��A�@V�m��֗�{���`�h���[�2�̼���	�8��1zNO��c;�vw�Y������}��[]AM��ub^�z"C��^�f�Xy1��|Ǹ?�7T�Z�"/��;����}}�J6d�aT� [T�X�2[���(�Gts�WO�V%a��j�l,�)���(��5��6��ݽ0(q�-�Yv£5Ž^���r�)��l��������]����e�.�=�e����ѧ�O����}��&d������u���ݍ����8s��d�����g��'��ӑ�-e�F��L�Hqf�xn6!����1!;�'㔢3�� G�Ї[���F�td���Dw�ճE�z����:��rH����gP�;��M�g�G	��X��ʖd17p9�Z׬���o9){5����K�G'i`��H5(�	���<��P�{��>�����ly��q����+��b�'��>	撥ysy	�lMf��T��:#��㮳|� p(�*4k��� e>�`B!��<�(����]Y}��C���J74�x�D�g��o�)y��V���޻H�F����
�7qM��kg�X�y������-w����C^Х#۝��Ff�"��J6�8�S�V�y�e�02�\n��WJ�̝�m���%E���槰���#��.,6��_)e'<8��$/�T��\�龊r@[ımݽ&�oT�������FB>&�)��j�8� ]�l=ҭ�&�#�I���cm��n�)�pp�<f��2��>G:R�(S�"F����~ ��t�P�aN�W�mAؓB��7Ⱥ�5���4���9��.�Hy�;�vrA�O�"Z�"�M-��������S�T��fE�A?.�2�e׈�l�شs��D�'aj�T�^�!#z��p@�&3�d���\�!cEM����{�I~���u�	[,���,u{�*��\]�#�G�� +J�
cdm'<��֋2��Ά��փ�2�;5W���G֓�}�+Zo8*�.����F�G>�16E�@�\KB�)6݋(�A���dG�}B��@%^5`]o�LѶ�������=_���"����16�gd�q�`�*����_�55qR��$��-�SS�kO,���a}A�����`����:D�ކ�z`��$&j�bT��OH��?W�C�y�é��<}���$�����q���s�T�����~d��+�� ��{I,f�F�(�&tX�y�F,o�,�O&��+i)���E?�T����k��dC*����Ptb�9"R�w��R�pz9O�"�b�8���p��HX�ŗ�ѵr]`y�|T���Q�!o5VvТ�0IF�]4#ZG�Y]b���4�U��eq��K�2���;�0{G�m�q����k�9ɿ{�5�/��3S�֗9-�����	���u���.g.h�Y"�U��w��Y���Zn	$w�
 %(�k�߫Y��n[r�MmGd��-��|�\$/��HG��ۥ:<���hA���G_���ғ�PI��Ca�C�y�7�[}7���Kg� p�n~�K�����	��H�ՃɅnu��`h.�L��_
�\�ߛ���={���+% ���f�� u�D5����RVWN/�3x�վF�L^���}3<��v��A^��,_�:��k�P1F�U��x��7!|\Zt۫i���#x:�-�R�d0�dM��b	���}x�w6w*�b��7x��EHw���
�*q=ˏ����c�^c��V- ����R�jiz�\2=�P�3�������XЋ�*}�Ѳ��M�����j�Q�Ҵh�_�b�{��b�(�[-������Dp�?�X~���HZ��.Z��Cr�R�3,�&
�a�Ris��h�]�m�����i��^�C�P��%V��ڊb���~ԩ"��A����������=ʯJ���{��e��� ���"+��&c�jQ��4����T?�������4��@�(8.�y�dY�.��j��q2T�:(� 2cc��"��C
3���P.oz_3�Ȯ���,��横'�&��`���s��XA��PfL�ݒ`�A���~:1�>���uNS�g�=*�%�$�6�x#���쁕Q�
.�(�#l�kT#7D