XlxV64EB    47da    1270(��\ ����F�t:$i�i0N��WRݔG=��m[����m����{�J��O�)"J�ñ�5��Ӯ��Y���u�Ε:����Xۣ,��|�,*�;諜��A��ч7��¸��f�F�ņ�' T�y���,�(F͈7��ؘ屪1	x�H?��D�"8��W�ǩ����F(=#P�k޽��<��J�{x'��q�n���sD�b ���Q�~��Ό^W�𭚐Z�T��@kDd';A�FP�K���>���f$��"@���e��e�oz(�����샬��T���)?z���䱢�,��ϯ�-fTi�hz�[�4�oq������8C/�b���0Ĵ��R�{�5�yv��ǖKe�����实��oaV�a�F��^�|W�����}��D�l��
;���s+U��&d{�!90l72���P��lH�m�_v� ~̷�$���]��ԘԷ+@�Ɠ|�A���Z��	�(�#NJ��m���*��T:���(��J!�@�'�Q�e1��;I�:��]A�����6u�d>Wk]��c��������j\,�}H4Cv�h
 �L�/bJp�o�����V���;���\�!��>��1�� �C�'u�Ǳ)?��9?c83Е�SͰ�O�;ū40w�A?J��k#O�e�u�U8�[Z%�ڄ2K�����q���@�bTm�q�����������-9�	�sh�Ҩ��nr��DScn�P�dV1��xd��5�vq�na��N�w��h�8V�W��]����4M:��l]��˥� .�u����Ӻ�O��K��$%+D�]aV�����JY�ُ	��Z�@�H59�Z��k�T�R����{�����Z֍�	��ƕG�-�Ϥ����Z\���<���0jk��i��1��C���0�_��|?�EfY֐Ů���@�
c�O�͋�e�f�"CJ����M��έץ���f�lDeB������=��&��5��� M,(۴W��tC,�dg�K���%>���C�	�{cMڱ��֛S�A�ݸ/��C �CV����������-'
����͛��w:�?�����N��fj���k=���۲���'��늾�)3����Ӻ�%�
	8`z�r6� ueWAə�di �1�?�⻼�kd\��(�4|��#�M���D��Wk=��R�/�M�f@iو߲�R�!ao�� ��`J� {��-��+h6,�u"q݅.?O&�Kؤ*���TkV:^0�[8Ryd��)x���"�-�0�S��NMN����~���(I�W�k�/,�R֜��ʰ&g�����$�՝�����L�G9_���&�n-o�3�-e�q��׼��V�?�8_Of�[4`K1 ( ��K��8���ALd��KJ�����gH�SZ�;w/�Tt�`�!a���1n����4<.��o�s�8P��8��b�p<���+z�	0��88�,���E��.�Ϟ�o�>�^����'�"� O8��\�������D<Mh�s��"ڕ�g�Oふ6�VY���j��ew2�5F�u���~�����cxU�S}�'Q`i�I��[J�U�0�Ū©������x+
(	���WW�B�؈<������ˮ�Wi�����C�k�d���Mf��0Ϗ��Q ,s��n/��tXߩ�/��!��QAX����}�t<�b�����8����y�"E�	�=Z�w�2��7���JC�À���ڥ~��؁
!�^���1��=
���(lq�V��3J�a�ǼU
!/�PV���`ϧT�(B����Y�\q���K��?
��yӣ[X����9�� �9
:H^6Q�c�&?�B�e���L�!����q�=��t)��:�5�0(���z�����f�5�X��8K}�~���(���:�b^�%��Q�m�*�12���\*�@0���4#��?��Aq#������_�Eۛ�X�T|M||ȥ��/��F%��m!A��� Ǟm�V����?��8�*;j-<����_ �S���*�?�xd{v�P�B� P��eJ�uY�ݐ4�#�����������Յ��O�!��7����B��o�(u��kV~��S�z4��I��:�� ��Lsb¢�lG�>�$t�n�y�&���������P[��a-�Q��`��,[Ŗ�tI�����0�vH<���鲫h��!o��Pc��e����p-�d�Z[P�6�?���;U�ؘg�^%m
/��e,/�`J�mWqI�xح�fyU�Ս�0O�60/A
����t	= ��@�9Z<�ek�� W�q��o�0=�������Eh";��K�@�l���&��������Y��s>@�u���,)��p�_�q���7i��`��z��-I���<�4��hFH�_GL�����2�7��d�d����6z�v���H�/Ru4��G<�;�ĩ �fe�3.�ޟv���M�yw��^D�-�9U%�!Z]e��\��NT�K��\�XR[���=ѐ�CH5{Un)���8���\%mo4�Ԁ�i�؛Z�j��sM#�o���\<�����d$���&��9e{]����@j~i���g|T� !�<E���3��1���~i�)���X�\kX5��|�#�7�X,��֟�g3�\,���iR�^$dt�(7�];��y�רh�CT0w�4�:e���׈Bxt�x^V:ՙ��* $F�S��W��` [��z�1kw�2'~J3��T�	�@�W�Ͱ�o>M]Ŕ�N����[��|i�6�b�-RX2�ܞQ�18�qWik��t#уn�RyÐ_�=Ts�R���&�7��w�z7V�OjGm�y�d�Qc)�}�Fڟ��=���	�·�h:"��A[j#����Nfڣ6 l*<���5��n�u�V
v�;(�bіN8E��-!�2w�{��j�J�}�,�p6����VJN��j�J-���������k�@��S��@�|^@�N�,�Ml������,��?��#SE���]Sۻ9�%�C�|PZ���G<���E���l�����ﷻ/���#�na���rm�$�p����Ĕ�V�f�gN$rv���8FWˣ�E���)fI��9�u�w�zw�L��䁃��CHwLǌ&_�5�t�V��H�6kT�
��{C�`�]g��+():�
����U�l�o9z��~�<,�_�Za�(3ʱ���B����,JrOf<� mh�C���H<�į�"���Q���	��N�m��#�` ����h��EfZ�p{�i9�$�-E/��Hr36�U[0�Tz�N�vۼ ��B��G��mj���F���^!�ՠ�H����R���.v��������x	��՝�~WA,kN�O�ĳ���	&����~.~a�V���A�]`���X�m�8q8�Q6��P+yjB��q¦z^êa�<�a�3:�S��E�l��y|<�+n��w�����8˂�|=
�����j�FW*F����qǻ7�3,l8�_6��{-Ӂuo�]
iV��$�]f\8ӧR4طZ���|�i�{S|w�=TI���8cd������0��KS�n�z��Rx L�ݨ��lٶ�W:bq�'1/[&t�g�4ܜ@#��X�O8����vu�hǮ�L*��-C֞;�C}�{s�˒�u&�~G#9Iby�ߤ6��J�8AMBIЅ�;�
���_��w�$�����^�e�kz�E�����JS�h4��b��4"��C��Q�J�����Rz��xf���Hiq�k�����E�u/n��f�:��d@r$~V �@P�+qw��x\��1ٕ���^8��;:��#BA�����.��Y��rſ��� g�A`G�{
I@$n[�"g��/�qɉ��М�a���<PXf�7��O.���z#F�W�^>M���L�����R�*����2�e�&���I�U�^�fdMla�D���B�y�_<�"���I���P�#�k�L��,w`+2W	��<ޖ�I�QVƏ�D�A����:&��8�ji���xVʪ܇d���c�oA'��K���������Ǣ��3-�+�Qs�+[��8�`a��C|�x�n\����V�/Z�B7Q\�r[�?�����[3���ߦ��#��x�VL���o���^�ŉ�n�D��>κ���GR����ryH�9{�r�	��������.X^+�c�;9�����6�(��
屢�����cX��X`��"bC�|��F|:��`L�.n.Y��A.Gsd������Y�@l��c|�?��EnJ�u:$0��C:�,�d�>���x�ܝ�X�˦�^ҋ�G�R�#�p:��Q����rg�r^�|�w!ó�A���YF�U�7��7�#�Eq���G�b��D��Ȃ�z��ɸ)�f�k�#�!$�1#�WP���!���f�m���Aݑ��BcuPé�8�"u�_�6��Lc��;�I�$�&հ��ѩ��+~��t����J� ;Ӗz�z���>6���9J
3{�}����2��t�R#���������z;z���	���k�F�-�t��x�8~����Lװ�L�Vl�B��%�L ��T����:@a�sM��ѓ���E���Q����Cğt��i��7d:NN�U��U�g��:�G��