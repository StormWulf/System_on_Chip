XlxV64EB    17dd     9a0f|!���v��h�����az �i6,�N͇��ё�t�yǍ�珖fЏ
ϰ@F�2�)��� `��Ж�L��
쾕�n�c}�m����F��mɯ��N�̶���5/�Q�����/���!���*���jy]��K�,ҷ���^��ɵR��WV����"��O�k��#��٩b��w賄�`�|�z��%���>4�XD�����%� �I�ރ�-��ң�y��U�b5����\�k�b��מ�;�2>q�9����y�旆����ӵ^5p�%�4;�&م�"�rX��?k�p^�B��aR����Z���׻�TCl��5�^��B�%��\C�)��]D�^��SxP�.�9�������zX\�f���ɟ�p��u���+�QV��l� I[Rܤ�zF��N�D�����:4�h�e��X�����=��19�"��b�f�r�*G�ZEL���������i��-�WCsU첫��1�����>D�?������>X��k�o��W�{�c�����z[�+|hKv��5����f����UU�ѭ B�A��)�Ax& �k4�RC�z!��"@Kh�=����*�|ڲ�Jj��M/��FR$�����{���F�*���gQ�	D�a>�]Ј�щ4�F-��dƐ*Z-h��:]=0��,��9G�A^w��Wh��-ozx��7�����O��$�?�`���뼹>������Gp���d��5��+C����R�.T�ׂ��N��⪅��>��&)���M���ca�*!O�uN�C�D�D7	��|h��,��sxa�5�7f��g�횰!q!��ˀh�ERR�{��0~�X
�~��{h��sD{I��W�R���R[��n*����{Fi�y���������z��&tJ~�e^�A�D%�t���qD�TRĐ�̩-�	�76��|W�;��;�������z �6Ro�ߋ���g��B����6ZN�rk�|���>횗!|͵�̂Ta���}�E:UL$3�nн1�B&n�(vy��:wR��L\ED��:&"A����&n����gr��HHw���ݎ��R��U�:�I�`Bڵ��#i�5_h�Z���h=>��#��ݱ��)�����ہ��on�7�<;����=��nꎎl�*M��?���9Y������׍���L*�j���$+�u���_e:�|1*<�M]����,����)��V��L fH^8�dƃ�>���M_��08�7����ccw�Čʴj�B]����*��D��=�w��b�m��yS0���v�7�u2��3 s��"�?��(ق��g��=`[�Ү����T�<3���U�D<��ܰ"�NU��N]&}�	D��]��4Lw��nZԛ���Cg�
A��s��&�}1Ѻr��u�z����=�=Q��'��fQ�յ4ɴ����?���m���b��V[c��W�~���U!�M�і7�}� {0bYE���V��^Q}���B֡~�RΖm:lR�ݖo&���*��K����H=[A�ge�e����O�q�uBd��,�����W���E4dy$o��\�&7��`矷 ڌQ)|��K���l"��`],�x��< �a���[){9�lngB�A@6B�o�!B�Ƈ��S����P��KY��U[^8�i5R� ��""�GS�Y��r�����wֶ��Y����=�,����h\�P�;�����Y�f��*[6?�mR��'�m��<z��Ѧu'�{661-��8���dx��_�Ha5�<p���{�eNs�Y�!��I ���'�q��m�����������!A��e�����[���I�ˋ�N���f�;(��v�[aq�a�t�~X��������*5�Y��c�.���!H�Z�B���D���h8��^^����Ȓ$s��[��+���"ik�mA��F�53�T��xe^��d�o?�D�O������p��%�Lb�t�͂� )���f;��K�S�42����:���x{�V',�5�4[�����=:CkԘ�6��r�S!���\H�����  �-x�������RDc@&���ΑK<(�b�Z�H��7�C�ȨZ*�qp(9N6�\ؐJ�@�:{��Tg��3ӈ���'w�⹼xN>]�������{B~^�4r�u�`]�]*���R��;N�����Ⱥ�]/�
ZE(�pc�@:��I�ż�{�:?�jk	Q&�!�����P�L�5ά�dr2�a+��B�6���KS��Ƹ�[k��xIg"
dz�H��`X���kƅP��� 2������1Po'F3@?v
�HJ߁9�ik��aԼu���s�sH/���i'Ǿ�����T��\��%[_��s�