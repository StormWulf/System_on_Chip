XlxV64EB    3816     fb0m�Lvf������z�3�ft����._�!/���v����V�4�Tx��Y�Cyq����P�r�IÓ��"�lN��R`���Lw�^��H��E��֮��]�2&���;c��ʀ�ډ���b"�1�|��VC^����1��F�e�.'A�Ӟ�լ[ROJ��`�ռ). jc��^��@��6��d����>�j1x4�N[���Y��_@��b�0�]d5��m�n���Z(9�'z(���1	�*�e�l$J�/�|b�n$����,t�<�iD���3�dG���@�R2����$�C�VNH*4WM�?��J�D��	i�%�a�	�q1�p�MMb�0~��@��0P[7ӓ�-vޖc	~Bɷ�AՉ��׾�b�\��LM
Gm馊�Im<ϭ˧�#m�<��b�:��4��4F�t�T��tt�bB#�F~�uw{��F�l�l�lkqd��6�M�PUb�:P��0ʫt�߃W��5���31+s
e�}W�̷��'fb�����O��V/����3եH�J	�)??�]+;2��kONA3�,2��U-Xd ����?�bO����?�wӓ%����wm����� � �2:Yr���%�/}�Rz���D�ew.�<�Z���՟=O`�����!*P�F� ���5�_��Y�jX��m�i?֡<xG��|d�3tQ�����MK�$QD������uZ��$���s)��A��ҧ�(CX�bG��ء4�N��:�0���|t�<�R����?E�D���)��'%j�҈e7��3�Y��X��'�d� Z��5�~C�%`B��=��AF�U[~&&���(��~1P�i��VG$�h��{ڰ՛�G��\u/5]�A��{�������ׁ��ls�O�4D����E�ԞjY�����:�o���	����Fo�����Hk�8��V[g��_��W�W��l%���i8�x�a1�dn8�D�K�T���LJ�f�����r�'WJ��	Oo� j��|�+�Z�5E������8��j�w0�h���{\;�M�^S�J��p������ԍ�=�����J���ѵƺ~J��a7��<d;'ܹ))wi�A��;B$`T	���	)��2�d�uI��w�.H�-��y��_w��u���U�Ȝ�Q�UI¶�6�m
}9I���4��~���3�ذ
	�3��e_C����N�<oF�a�Pa�I�G:��@�ǌ�Ά!/�~��2�ZW���!���I�Z���e<r*���4����w�C��U<:�f�m�E�ߺѢ�O5�H�@W��f���'�y�7��Ll�N<8�f8]��b=S�����eDd�H�[������d��K��q����u:�xOR��gM�D�b_�/�L� de)�I9J������Jqq) .�k�?�F�g�r�r��r���ȥo�z��=`�9�R���+���:$M��Խr��,.xir{+�iGRC�����Jh^�q��L�cU����_+�X�+{[�cp���ڣ�ʑ�sO�<���܋"S��=�Ը�1��7, �3ƾ�Ρ�X����sv���P��x�ߒ|*�P�nX.?ˊ�q0�6��[�!\�Z�1�J������ bl�.0h��Rt����S'���/�����(8���i�H�O�@���^f��N�pP洛|Fv��|��3���(z����J+�O�sE
G���2X��Ŏ=9�:�Ɓ�`�2r@����U(�/
�8l1E����\Y�>�ZGZ��,��S�\�=��R<P&?s�@9tv���cG9�x � �@&��ǅ�*:F�J����K�sw~�j�3)GF��M�OX/��y~�	�s���bJL'^���9���ǚ6��$-|�_E��6��Ԙ,�"���ꨈ���:x�qb�tK�E	�s���|{�������8�>�yl*��A71����
!�}��:5�}%������UJ����0��V�d���!g6�O��3F�\��k�X�<�t��Ñ���[T�^E�iyF3����gV�Q������d���s{��jRq���y��t$�.��
n��嶗)Z��2��&�V��tO�{�i�c�J� �SsOv�S��;�#��R'��s~��y)�ֆg?�<i�]& iPNb(��I���&�f��\� *��&ҹ=)���{�G��ڕ�p��6�%k��j��I|g�0�8MVz;�e��B[����eN�ۅŨ��z9 ��۲g��n��n~�p!��Z
�4�Z��Nq��}+�5S�pd�ˇ�������Һ�����93��`K�\UwP�>�������ē��^�4�GHj������m�!\P�!~�׸  5�Ȥ6J��'��bi�����[���_�d��1Z*3(��y�N���C�3����`�i�ϣD���[VE��[6Ʊ���7����73�9H_�F���k�Jh�f�E?�H�Ū���e�mƈ��Bt�@?	��<�5�R��E���
#[F��'�k $Pc��m���㋉�i^C�q���+o�#� )a��E�'L�oi����Z�hsӞj#P����?]E
��(�	������?�f���lm�����W���x����7���F�rH��ظ!!�k-���œ�il�>�ѻk���f���Ë���V�>zCҧu<Q���Ū%}�/�c���'�b�r��<1���<���Mq��u���'G-���z�1� N�j���Đx�"8�{������^|I��h���K��G5�|���ɗ9�4���#��9M����FQ�d9�+[y���7���ێ���5�i��*�d~�{�b�RYh����b �+?�˪���Sm�(B�K ����M2j���D�ڪ�k-�B~
Ւe�Ҙ���+���5�[M� %;#��3vI2|�'le��~gmh߈��,�Թ��9`�)ޔK��?�V��X?��`tf��b�؊$!�u�%?�d11�����&8�M��fs�?&��\��na���ׄJ����zkyM��>��;����M�����Հ�� Lx��R+H�At��1�O�X;��JO8/��"ƢE���dlE
���w6;@%~��O#�VK��;��Τ�!S{G^Å�i�ޛ�;x�C2u����������m�,w�j�7��oQ�W�)�H�ձ"��clt�p�[(�"� ?S�G����O�E<_��w�evcg�oZ/���iV:��ƈx�~S�Cum����r�;V�ƈڦN�H�ZS��S��<�خj�#�����	��/�)��!�j��{�,���X���S���h�60W��-�˭�/�?���n!�3,&��;�2KI�Ӽ}Dݟ�Cλ�f@6�ޮ{DIN~;є6%/�(jq�M�����:��Gc=�YO���${����c��f��fyg���,!ўZi�>��z�E�R䦃D��I����@�z.o �T�4&��8�1F�"�YQi�@D�sS���,+���x�� �	i�r��9W`j0^v�:Zo���łn5����wm2܇`�u��y� UT�Cf��Yk��S�eX���ιv�'��ð�D�-lu�w����i��8�r	k�،WM�����TT.���E=�ʭ�*.�٫�e�A"j>n�=�Ņ���H�s=� �~�B{��)Ql'[|w��V=by�����=�wB8/IG�����@��21���ƽT�}��z���#x��$��R᪆�� %]��{�V�]��Wf��E�={l(+Y�ǐ@�Xh��;���}�:"��ST���n[��/�}h���z�S�X ,i7�/�9��!G|��d�6G)mOZ v�"y[�oPO�_�*��+*rNz�����䏚5���0I��a�bͿB]ݜ�Eq����MaQ�J!