XlxV64EB    8541    1810��$��T.�>�7�Ö  ��ց�����x�� �!0�B��vxWܸ�׃	�z�W|!D�D[�
� ��A>�m4d����#����_���p�U��[���[K��P��T�.3�X$m���Z�/=z6U�39�.λ���v|�52�P����F�C��no������&<em�h���뇗$-=K()����
�(�\b���f�U�ޯ�ˤuG�5���B��Qv}D�����Vq�'��25$�"Ց:�_q�Grx�<���f�wm��2��X�V��)i֌1્���R�W���('��A����\�ˣ�1 !2b���z��aeF;��oF�*��jC��cD�Q���t���}p��4~�e2�-6�q��ʯ�p�9Z��2��%~���+��I�u�9�sm�P{rp,�9;�:X��!:�c|�Z�晉��jv��'sRҢ��I�&)�l淟��P�Ѹ��G����������	����F�+!=o�۬�Hp��o�-+e��usv�B������M/��^��Pp�0b]���;v"�e��5,�p�T�$���@p�]����w����I�*�5�]��*F�^�b�f�E���� ��� ���IK*��	����4���y�UL�|�㱯(�1���T���k~�.������l�!�Q�
ܧ��A�q�{c'����~��4�JtoJ�Cvk������6�*'�ڙ�Rl�X���=���CYY�o���$��|���؛buu���=�"�z؊S�_��} -���H�<��*��/�4|p���L��#:���k5%���
rv3�����CR�VŚ�}�7��E/ �v��"E{�?�8g}��`D��%�8����9�cgS1�>��'�No���)�/����!#�Xɬ��T8
�qlb�%k�A�;8w���7��n��cШ$�[��d�/�X�ȁB�pTdd0��z��S�w����c�)]�0�^,��s�;%<J�����E�0B�~5,�5m��-t8c3��>��f����a�Wv�$,�sdl
�»` ��=u��=C2͍�o:^垖d#{P�h��	�v\De�Sh:��1Ey�z�U��R�}S����g8�E�e�jbZo�`���iV�ˬR�'7��"C>i������ƴ���it�)�����+�}�&=8�~F+�v���
Oq��
�Z��7�ٱ�̢tN���L`+��/����bb�����m=���OT� �@�Ɯ�O�_�Yӆ��e��C�g��.�]1;���kI>�WR�PrJ�?0�]��j�{~�-*y;}A���w�~�ʭ��\�Y�V�ё�� ��zm���?�*�j�\9z��������p��Oϸ0��Gb�]����pE�V}k̟��7��WP�v @�������Β�1LC�T
ģ��F�!�)�#2��2~���+��/�^A����aƲ{����W�{~SH���iu�@�"�v�0�D=�g^X%��D�3��F�yO���x[P
�lȕ�����b�t�BtE�^!g���kh�]DY~���#��$�X�|u
_k�Y�a��5b��a���\��R�$�A�漉�K������\���!lێ���9B���J��Ly`�� D,Z\sM6�t��إ�(@����w	$\x4FaM�����S��[Cf�Ơ@��o\�ܳyt�Hi��d��p�<	B*�����:$x�_�:�Z�D�z
B�i��RW��6��t5�a$J�z�k>l8�j��a�"�|z��7�����xtT���R�Sc�:��%NX���Jвa�4�i<�8�*西������=Kj��K6��g*'7�e!��=C8��_�Nf(XV;Ъ,B�ϔ�U�BVQ�1��KX�Z�x�8���*��|�wAj���쓏�L�{�Ƃ,�rH㧱NO�y=w�'�Z!��ُN՗>ٮc/���\��T\�:kT�1Y�U�>�B64p4�\��FM�� \���}���d�1��<�ځ9�yoo`(�-|&u��&��WJ��ҾӰ����Z�H�0��?O �` .�{�W�����O/T�� ~��h����P��x�Bp�C,a�����m���E�$�u�#  ߼��}����!QμA6I�aU�_B-�=B�^�`�������n]!��<��u	�5�\�יִ3���\�(`����S�� �� �Ov�	d2�^��q�?�Ĳ��;��_��qwt�7���ˈW���枌��Fk^?l[?�x���"0R2�M��b��R�z�-����Yϰ��-��/B݆�d���.t�|a�l~J(?�S�
���bo^\�E�k}s�?�%9~��1!ܨ�q����l#���l�O/��!�&swݾSR]l�4�݆��ގ�a	�ׇ%jΝ���ϟ��I���n}���S�i�5�aP����/wWg��e�N:� �Vy�Lb��=(k���GR��M&8w0�%H�0�^��I����,Y?6�T_\�����
B:L�$�)��f����X��Y�u��E�!�ÿ���v�\���5[J��/���r�&ֈB~��|.O�}ī�pፄe�ݽDg�%��Cn�P׷�T% �	���k'�0Y���XHi[���!E�kN�K�X�Gʣ8Й�k��8'��ơ�c��@��w%���x��q�{F���R���w�8>kD=���t�g�4{T�,�Z���=9����B(��L�Qz�w������aicI�ֲ�]J""���9��H����&$��]0z.Y�ɷ��	�g��PN̿|��,m	J�T�ڌ�Ѕ&��5�d��Slh}3���ݭ�X�ZK���´KtUg��(ɽp*]K�:�i������L'z���Ӕ��/β�{d,J��a��`|3V.�>�Na��zB�H�7�.�������k���VY�N�'��26��)ߣ	���̎��_�Z�E��Yga�F�g���!P�l�aK[o����hȺ�d��yv�E�Ζ�����fɐz���?q��.F]*���pc�����y������W�;����{x�S`E���1�!�+7{-P���۾GIp�͌����X��}�6l��}��:l��/m��}��0#���#lHV �&
w,Եb�U���,�?
�q�<Y�Ԁ?RX313�J����9UmcL�H�Y �܆qmm�R��J}m�}�']���G}���.nA����4^~�w�a�&TF�Jj�c9o;�$[b`4�����I�i]�B�����m�ؚ����u��8�}�Ō����Xب��`z���Ń�v����v̗-��Q�M���l?.ـO�ٲ�N�R��H����N�NxfO���p�B��²�E���d����<Nl&�� #ۂ�v��a��y�kp��j���H�a��X�*v�1"��;wD�pp�i7�1���p�szB3��\�.�R����=��0u��G	::IE{l ̺�8�|Z)�����DR�f�ɒw}�_�Ɗ���
�>Y!�9Z:�x1�f����}�ʮ����`J@��3�����$'�@�`��ВV��� ���H���D4���ɵ�Q�����PA����j�1S"0�bA�F��e��G�đ�& M&.��d���&f�S�_��MT�H/�ّ}��(Pq:�_�m	ȷQʝr_�h�&���)�	��Gb���Imc=��3�k�Oٙ6$���ɩ���q5�,ta�?6|�5�ʭ�3����R��6��J?IQ�D߬>H�%�%����˄+ n"A�v�!���W=/���Tr�@�=��d�)�#�FY4�XF}Ho#<�����א�q���L�L(w I��a�]�)���h��ի%9*H@zK����0):�oi}Kv�6NQ��i���
��TNKq��Kmŕ�e�]pR"�\��^[N;b���8�I�m��[y����z�
wK6S����}��!w�8MG��9���`>�Y))��N�>x�_?���� w�wO���3���;��ԡ��� �� Ȫ���q�<�	\("�d>�*��G4��s���#��S�#�_�{�Xe�J��M�6\
'i�G���'��Kz�q��?P��*�o�"̨.�9%A+/��rF��I�On��$��	q]��'���W�I���fwm�ͯ�;��g�e����F�@���b/�h�.��Rݷ}+���@�RHz܅�/�d|�o�`O�Z}Gȱ�C���w&%//$	40��%�՛RI}5�dq��G���U�ˌ�2dcA3���%㗙��X�:�_*7�;���Eq�v�xm�,���|T��_�Ý�V�u\�)�;��E�!.�;������!B���
d~�<�b�t~^�T�ʟv�f=�WY��H�N���$�|����Ӆ�~(��<�C�/m:� Ų������*��֤�����<�����|�.gsc��GN!��Z�ə�p�X%
�x�c$���!Zb^]eK-�_�-M����%��)~�竷T�p�y�a��}n��2[�ֽE��q�a�Yo.֮sBuh�Nķ����#`z �wQa??}!ɚ�c"���y�N����x7m�^���tI�1�K�I��B;c�y���d��`��ё��z�Y<�z&<��A�7&���o���:g��^hO�{G�.�01�K��#��oVr�|O�ν�e5UW(�Q���i�>�ωGa�`+�1>��5<&��{$��@>��ڰ��ӪΨ
�g�2<׽²�Gn��?����(�Θ����ݥ1��e����I�/����� 	R��p���ɶC�֙E�+@��@O�J"�d���|��ڪ�G
��Y"��/H��І�wڃ~�Z�(�F�O
�c�u	��@�+o�&�a��fc�I���l��OR�m'�f�щm�w���ԧ�Ή{� urx�z^��5&e�W� �<��(��Q?Y���^��R��������<C���F�i�˴.�m���߻�*!1�"W�D��n�PpO�Y�G>�@�muz߇~�/}3i�уlE������G��u�MȕA���)=���vq�SlP�c!�co�5�J�Q�r��(�	��U�ߪo��m(<�Z�� l���(-!l�Q[Uw({��s���W!j����X�vd��:?�k,%�j�@s7]"6����!���N�DS>p�8=��>u�X�-��Cq������A��T�i[�}T���@���E%�)�3�I���uE~����y	j[�6*ud
���Ii��^S��2]��1^���j���L�D�h� ����/	�o��M���Xো!B�g�(N�oz�.���̬�1;FWઓƃ��m'��s��Wf����4B� o��3��iӝ����ߡo*��#����o�� �#ĬT�Y'H5��4P�@��P�fNL�~��0�o�~٫S���N�URS~�7�N^�D�땈3Š�I<�o��TŌ��BpZ��l����*CP��{�/��\<�3�@.{�B�a���jqFZ(����i�E�=��8�I�5C� {�h1����]�
������ �2D��ϻ�oZ�#f19�c<�c�U�=�c�'�Sj�|}��8����%�/m�<��\o�� *�r��9|(��͎�b*nRƓCТY_6P��f�]d��Y[�)mOZ�>:���G�Bn��!��Q�������}�ޅ�]��T��o�ĭ�b����� �$�����l�p͝7j؜���R:�p����q�'nbCJXSJ��4�h=d�6G�%��h�ɷ#�[��/�����9�ٸ0F�
�p'�A>O��L��S���@�M�O�Z�V� @�mH)I}��G�>��r��4�;{Y��\����V	;����3q}�ճ'�����&!�ꌋ��{�X��ﲨ��Be({"O������<���M����w´R�B4)a6�65K���J��f!&Ϛx���Dm�R��.ۤf���^���OKU5_��2t�H���'Z&?rS0G$+���B��