XlxV64EB    431e    10b0�e�Rب��r7�Y�bq^vx�N�p5'ǹ�ڳ��7?���ɜU�|e\��@�����ZA;S\F�Ԡ�6���=�C+T��c{�?�p&�ٙrM���-�ї������sl	�MeF"��}fTV�;��;�ں2x��IeB�&t�s.�oz~�P�F�&JR�6(��-�� ��]� �zc"�_��/(�Y�Z�
����W������,�ee�Cv��)�}M���S8V=g]?M��@��\7;��8�N��M:����u���6Z�G;�<�\Pe�E��@��E-�z<F���v��{l���<�\E]K�X�]ka���c�y�����-�������MA���	�I����>h�[���^hJ2�PgA�u�$z�J������b���+P$F����~��{�&	 �Y.�(���5�C�������S��icSi|
0Q�Rत	�SGm���h�]
¶�o�Q����x�����g'^��2�1�`z�v{|�˞%�������H����r*��_��t�L���W����5��b�Uk�e&eܭ"��X�ɇca�rH�9$�w�����w6M|��q�ا8���+"�G�K�s�b	�nVW���jN0���oyE)Eך"$�������BD�K��'cvo�V�;0X�y/�@4�C�h���w���e�>gO䭌s��-���?�-��(���M/�+��� ��]��"�)�|U�Tx����%�T]|�5T��|�{d���M��U'<./��Ʀ�--�7{���#Db�k�&�ߠ��/�#��D�d+�P����S2�����Q;G(!�T^���X�I�g��Z�ޡ��3�����9DC�]�(�n���01\Ǭ6ȼW&)�����}�)QϹk/�6H}�h�g{K}6e�����_��2\�x�S�L9��9�Osa��1�������iVksX@ ���M�3��3(A�q���ň���ٴ���n�~i.ŕ�oW�{�O.�nw���O��%5S�d�������X�ǫ	�W店1b?�֗!n~�qgɵ�Mx���6�]��D�k��
�'bWQ���ɰ�؞���^�T)��re!����Q��mjX}q�*KU7�0iJ
���
�[���R�(�#Q��2ƝM���/����c<'�m�*
�'�j�2���גҲr^��e���.�ʰ���|{�/t�o��U�YʕbhUmEF5�q
�=^P&N<��2�O?\Ik��A$���8O�0I�
�uK�Ȧ�4��9_�T��'N&ʗ�Ƌ��|؊L�D���
�N��%D`�f�eک����6O��i4J�/&�Q,'vxqE{�@$f�0;0v�[����8+*�,,�8���%���"1�Jk�,��}*���.x���x��s�lk])	�n\;|H:�j<���L(H��7GM[@H�9+mvO����ؽ.��a�u|���Ո{��^�<�b}5	0���J#�ԫM����"E��P.�eB�+Y7x �����/ꔢq����3u�K��@�`m�(��j�I����i�|�k�nK��0���z��?3��6x�5X���w?�J��s�{u�@`u�%��I1TL�}���y���M�m6
2���c&�d��g��[ލ7��/)�f��C�QLzb���PEN20kX��~_���B-a*+f��������]''ﯴ޶`���"�\ԅN1�U�# :t��� ���l��	�=��k��� �qa���`|<�eM��)�Z���m9�
�펡�\���[]B�e�'(���y*F��M�V��i��>iA��%�K	h���3^h;�q�J�t�+OL�dB���hL�7txɴuk�c�Mb�d��]�U�A1k�b�7
�s����l�AD�	�Hr/4y��WT���(�������=-���n���).vT�.��Ӱ`0����w��9�>�s�+�e�$�������4x_=$e{�1B�1�㿙�i����X�O;7Y3ɷ �V|;.�&5��u�d����irGlk�j�����Ml�Y?P��g��{�(R�@��B��C�7C�|��R�N��YU��)e�{��oѱ��;b^�\��;�"4��V��J�I�N�S%J3{���y��.�ʞWz�3TyZt�t-�c��`�o!�M>�^�s��*�P[�0cfQ��Os�Y҆	��2�Α�xPh�����!""�/!{�u��ⶰ�� tڝ�5Jˌ��<!�.o�>���$&���:��B�k٨ڪ�&)���������/K#��.����!��f2��"��#P�����]��k�=���i������zR��c�g��'��]2g\���/�mo���X]�
��v��َT�R�~6�v�6F{��f�Ƚ�f������Gl�_ҽmV��5�×s*�� 򄽶QS� )ud3W���t&��O����Ē�/)҃!��&H�3ݮ��J}�{g����`e��ܙV���1b:�=�^F���h!r9�"d���]���ֹ"���3�^���Ī�:�?=��L�M�Ʋƶ�V�$T�q��)�S���~@å���5*5��K���*|����:+��^��k[�Yby����kJ���R�~��`PՔI57���>z��ô~*q7�[���ߵ+��r�����i~����,eg���o����^�c&E��Qb�t�.�V%�ωr�z[��6��9#r���%�l1��M�i�T�z�����-*-��?����%�k��2"�fI�<�2�����?��"c(륱�e����Hhv�۽�(��:S��  �8O��\[ �Ҁ�l}�ͺ��X4���\�:L���^��"����9²觡@!�Vg�7ɸQ�a�bY��!Cw�}���W�wS8|ʤƦCu$�X�FH
8��`�:�7�}����ޥ&A�uLo=ĕ�=Ӂ�*a��¨2�oH�^�~ RzGR�(���� ����'[���d�E>���Db42���k�PM�ﶜ>W4���N�<*�A)%�1��`G��e�����T���JU�6��������]16b��A@��E�ABo��-�Oh̤t��"O��N�JG�_Z<A���\y�`�M�_�T���,Сy�F�V1T�Ng{ ڷg�
�lH�(Ve�g��]�ZF�Cy���4[�����Kk�u2�GC���{�_�~`t&�=6�
i$x��u ���}�=Q=���~�d�5���@H7U��,��$"��j�7"X�=�뼌0Y���:�>��@�1-�CL�Dǝ�1�7�;��H���;�{�~��qv)H��a�H�
Q�ES�����GGؓLj>���N,��6z2�}�v�xwTH4}��^�l��_�Ǣ+������ X�Kn%Ei�2����Aa$έ�9��iK1��Va���w�<,���]��
ْ���>���n�֘�sa�Y���v�ˊ`v����M�i)#��o�`ޟ_�e�N5T�w2�7+9A�p������u1���d4٥�+�$*}f�3�/�9���H�]Jr��) քg&,#C��c*�H�����n�OP0�4r+O͊J.lR�2�Q�'D/����,�\͡.�"FC8@��?��C߆�,�u�4e���򽋪��6{Bkmwx�{�!J
@���$HX'.���)�d{g�q� ��g�l[�ѭ�mgۉm�$a�=�O�R���#5�*��8Qn�v��Vx���!�Ѧ�Wa��\�IwT��<��ǯ�Od���R� �`�
pk��;O�<�y�od���450�sݨ�'bP� I�T!.)�'|��0.o����%�Ԁ|/Ȯ�cI�.�N�	#����K
h�/𘨄�����u�g1�E����;)0�B��^�帴�ͿO@��I�!+��,�>a�m*\�0�6f��^�
�n��U�(�aa����x�,l��7j�%��f���_�M�ĸsԺ
+�D��Hf��E�؞b�4���VB!�a��8=��g��3��IC�ڊ�?m�  �#�S?��R��Yj���0~em�xo�R �kJ�S=s�+L�J��.*/�q&�ܪ�����nU�N�4"^mD��$Dx��p~r�S+u9]�b�P���aU����E��M� 8ǭ_�w*��h��Ϋ܍ɫ��-4�֏_ȱԵ�Wp�Vz��op���t'�q8�u$\���