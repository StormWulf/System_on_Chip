XlxV64EB    fa00    1ea0�Y����
wU4]�I�_�6qX`�fK���;�I��Rӛq�������Y�v6K�c����pŐ p >D�qx�P��nXmz�&�!��bS����,B�r`Vgx���Ѵˍ�ؓ��6:�(��Įi�e�Zs��d];�D�MI�nK�#�Yi1�ddl��d��9dG�)Wˊ�	����&Z/�rRU�l���$# ��#
�4��!NeQ�LH}6�9!6d��?��~��K�ؓq9����vC�,���J���S�k�'�)w��+Z�݂��d��T
o}|�, (�~�d���ϴR����w��l?�CZIE4.*n�tE�D�l�[ٜ*��A[ru^uom�#��2�jTV�s���{�!) KY�$��y���-�OL�͠!K��$���o&����EM��3U����^X�l�G9��]����}���.c������'�S�Q�z���]ǅ�����f�~Ϲ��U���2��G��4���X�v�	�3w͝}>6�̵#�*n��t�R�@&���'�[#N�P�w��ȕ���|ILP��m\�
�ܑ�=�2��'G�8�� k���>��o�2�@�௏��$f�'��n��۩n1��8���e��s&>�Z���|qK�nژ/�f\��o�DV���0�T	F���ƻ�c�Ŷ=�lL����C�o��>�J��1oC���:��+����2���h�y�k�O�����j�J�R�) ��ǄK� �j��Oy�����W�pT���v���
��� 1�$����G9n��-R�^�ٴ�6��$Ã�xć*0G��qV�Zi�c��LY"za��Mg"7UܿW@���]aAy���8�Q7����)/H�Y��:�����.̉��^��Ց�6c
�' P��|TY^A�q��֡�����Wir�h�� �i�?eҞ"Ku�M�VA�<��@St�7H�*�Dy�����x��'�*�!����������Qn�@%���=�S8��	Dv�7�_|���>��ܺ����bH���|1�M��$\���o���i�	�0@T{3�FvB<����Z�xsH��H\kb�T�#*k���<�(ɻ�uɊ�oK�VÝ���Ѕ��A��,���&^�v����Cj�I�!�3%6�qt��nX}1���W_A6�!�oî��n���kɺ1mf�� 6N��� ����T:����P���S���BȠ���2$��������3��1x�ݵ�^�큁����?T�Z�4!i���ł?Z�����qe�FI���m����r�Io���������ŏ1|������	&%{E�QK�y���UːPbH�o��O�q��������C�sܮ]oJ��,���=O��i�����I����l!���V�8)���^f �������I_���� S����L����Ec�L˚D�t�+m �2�(�߁ÊH�Ō�g�#!�=���*k��[�����h�����5e@�����X���AT�Rq�.N���u��@/ML[y.�i�r�E��f}B��2L�ڱ�U>C#�Z-����xX[�fH���x�g�b�]��!+�*\��E�M��JI�_�Vto�7�����
��ʶ���z�,�6��d��έh]�MLr����Kd�r)��a�;*��E�B�^��r�B�<�>�v	�v7I[�v¿Ď���'���Q��'����W���=.6�%��K�m�R=�c��u|���e4)��ͭ��أ�I�v�M�ƣ��z�0@hO��y��z�m%�=�ݿ\����JßhAIBk�P�7Zh����\'(�?621�z�" >��RrTϣ�L�C��q�a�c��K�+�0J�E}���L"�*���i6d��i�����Y��v�����zw�\� �.s��)�);9��ޒ��)(�$��؈y�x ��,�%�����I!. �co�� �_ɕ�9	CC��p���}�*J�o��ł��U)$;am�iN9��cY�$��g�!�e��j�C���J˧+@�g����+���,fnWjɿ���営��6��.հ��H��dEvW�ؓ�3X����}�\�Իʽh���u����c.|��?M�P����9B������Z�p���f����1W�V��Q�Vr�"P���9�c�x�)����O�ܒ����^r�Ȩ)<��L���ߕ�����8�����T�uK>@��7������4���Dw�r����N�%d�O�c33#�g#.���N�ڹ�a�˥��Q.��7���ܴ���y�u��U(�ۃ��/�$�ʽH�ARa^�訄��`4�����6�a!�MG�w�V5�[+)�#׆ڬ�.��5�>!v%L�9�"�kt�2� �Wa�y> ���pp�U}-��h�̬˄�wV������#D��i�����7��4~�F+;(R���r�i�&����rWA.8=����p�g@5���]�O��o F� %��Nu!;��s�6�Z���Y�k������v�u�ۄ�5��6;I���R6T6E�ק�e"���(wKR����0E��t�[75�$ܥ>Q!_��<��;QN���4�m��t`�K`�j��W��uW���{��Ie��msŅ2]�0��k�'�#�u'&�8
d�d��oxڻ�'~,���\9�%˽�GGN<�0�ȋ�U��KBΏ���&��'Aaa�˹�W��µ+,�s&B�ﻪ��YͰ�t( )M
��V2p�U� ���Yה�=+\x�M��˦�?���@�+^��u�z�e��Z��B��S�pPTU"��.PN�oP�M�q�q�VHǬ3م�Xν1?�n�a{��ה1R27T�XWq�w܏��C�#f���Gd�K3ݘ>i�js3Q>��4b�)L�pD=�T��_<GR�R� v��Y�}xk*���Y��hox���bA(H��z#b���u1�!Ond���,Bh����.M�Ef�l�]*C������+OG��Y�@��m3+s̰�M�Z�=Gl���L����D�� .�`����]���EW-d)�t�S�"��P����^���¨z9�	�z#%���p����� �	�������_&x:�OÙ����0阻o�����u���bEI�ŘM"��M��j`�hj�	�w�'_gt����O&���[!ْm�o�Gu��hR��*I�?��桶ҁ������<HȻwu�}�������[8Tp��^У��Z����2�e��NoG�]31��&i:p8��G���N���,������	���tS�>��z�	4cH�b1�#�ڡepc�rS�}�y�w[l;�c�����L�:��=j�]XXt�G���&HV����C#�g"���
����tw��F�>�q(B`��#���S�{�H\ɠW�XeH��\a�4Gͥ��j�$X�ؓOy�"����G2��A���{o_V�|�r�	������y���N�F��=�i=63��ª>-�}P�0�[�G	�ֈ\�L+��F�����d�����:�$�"�N)�R�;"�*����6&H��媳�E-[�+�*_ڡ�&�Ãp*z��7�-��]
|@5h���s1STA0ؑ6��̙p��V6%�9BP�²鷚0����gH��e�f�ڌ��K�c�^(�~G�p�w|ҏ%���43H��]A��%��-M�<D�9X�5fz��&D��s�ӘR�^;��v.|<�ϴ"����l>0�xޣ!t�Ud��f��%�2�.�Ya}ͪm�HF���(�3��޽(�c���l��2Z��Hl�ah�~O��e���!�=���w_D��[TQ�̙)ԗsGW�*V�[��݌�\9��A��*XU�r�b���:��M.�����7�N�~���TJ=8�r�H�R��Ҝ��
e���ī|i�+W��&�Q�$�� e����e�Wf[ז6�?�CE�������e�2��0�����Q	^ł'����d�ڙ�����f|�����c�f��?�y0�f�n#��ci�	��]u|7�k/�d�g>⧁��~+W�E/j�1�f#�ǿ���ʡ�ə�0d2F��$�p��h������v�KoA��kR��]��@C��+,�0���X�/��wQ�~yQ�-�M�)8�_f~	O(Gh(��GӞ�e7O@r�9R�Pm��.��Cj<��o���������'��,c��d!|[��9��жm���.;G�w����Ē��
ݽ�,��[�Ծ�����tA� �`	3��c��<��!+4|�d���=A]���^�w]��q{�\�����P(�o��$�}R?���nx~|�а��4_�/�܍��������^���ͦ�b6G���Ľ	9ˉb�>dۧu��]��@�]ĵ!k�@4m�JZ�K澵��>�Fӝɽ��Ϟ�9�G���3Ȥ3݌�6�ҕ��K�����T��	�|Z� �b����#m8�V�a6�DJ�&�-���1�I<N+4��&5
H����7�\��u�1!�h3�)�F{���-�Ǟ9�m&���PD�h��F����U97Xy�8�+?���B	C቟�#�p��^|_�l, �d�\��;D>;�E�-�6W���E�C)�=tk�Mz��9���d��o��N��)�$����R�t�	h�5Ft�ui����~�'fVcv��S%BD/�m�k7�4{Yf��nP�7*�g���F��
�V��Z�Jl��1XY���=��m4�����!���1Ջ�I޻�F{��@iVvE[4�;�~���(�&��w���z��u�� 8�ǉ�u\*��s�SC�4&8��~�r���u����G�V�z�Υ��7��;��5�!'5��4���]�b��G$:AN�C�g��*w�<�{���.�4V*�N��9z������3Q����+��(�٬B��r�P��P��!��@f<���v�Q�/Mp`ւ������Q�A���~������-&$�K�����)�t}�,�R-[T{=>w���A[d�p����uFk�>�W±y�,�`���lj�tu��d����+XIY'���o���Ӗጦ(Sv��Հ�Vb�GX�P$�?�G����RB���-�s�d�����h�� ��������Tٰ/t�0���}H�Vm���,�{1�Tڢ�;�KxS��r:Ư����eƆ�M�8�%����E9&6��+�e`�gI�\�Ľ/�J�Xgá��m
na0��f��ᙓ]��*&���L.�W��� p�՗�/�WEY=�#'�|�\�Њ�zE�l�(��"�ԇ�E���.SҼY3��Q*�����������@�W���0(�,�ǖgm)6F��v�89�m�x�t���0tX�=�JG Τ3F�ݝfښ�Fz��
��B;��6�h5+7��<6Q	xDCT���Zۜ+�@ir�%��~[d�=E�4�^
&�����a��|~���A��b�+:����#L��	N�j��Õtx5���o٣�|��3h�4m�������O�)���AgTF�`EY��q�Ou¥*2r�/b�L�4�
�z��\�bS�z�҃v�+��,�IP�݊b8�J:z����ڧ�z-����F�z�P�Sb	��,j�u��f$�j�\�:/���~�sK�l�;��2�8-�g�F�a�~2��Z���Ȗ�y�5��U9>N�b���p�ύ�J��)��!�Yso��55�q!}Ck)�35>ҭJ6Y�YA���F2(�1Dt�p�x�eI+��ZC>��ȸ2_Y�x�
#h)��:e�|� �����[_MC��{b���'~��ĸ�Nk�7%[�)��h�ظ[�xܿ��/���O�߄j���2i;+�smrTqJ#ɱ�̞�sF�/yt�9ޙ]�C�K����<����ƣ8.�Qx�wB�{����}�&t���`*c�uc�OE�Ś�w>+���y�d|�@�e�F�:��Ɣª�,��)j�P�
˟.t�g�Q@�@I�;%}!�*gIi�9Q��>|t%�ST�53��@����־̧6�GE+Ie�?3��/�Y못�{;XT��C�6��m�=�3X��e�D�5Ǧ���zZ@}BVl�����#�#(�Æ|S�2���C�y�Qa�|8�����6z�e�:lv'���SRU/69�-� ���s.բ*��`Z]�5��+�شuκ �؜��͛/,��Z�W��Һ����h"a���v|hr��I���W���+�Ū��o����z�Fs�׮�p����<E���V�,������1���忚%:�y��ĺ����\K&�m1���X{AEm�G~"ǐg%�#Y�񏭄rÆ�d�|��yn��V����4B��f��S�2�����̽ul���M���S����p}�A��+�2���-C��� �D,o��̀��O!�G��a龛! !P��t�(I��O��O�Ui����B�*Zh�G���^�ܳaR�jM��Ypn����Dp���?C�Ǽ4foCE�S�M�n.�!�!A�%���&�~G7K	\�i�rA�P�#<�^W�F���jե2�m�ی�ll�;�@�O�(@cu�i�a�wmG>,p�I	Z�v��cr\��d�A��=�mO�%0�n�"���g��S��,8ΐ�y~5)�B�%�N�e��d8e%�v����U��mT����M~�� ��b�ee��r���QyƯ@O�ޝ*@m'��=�,��mѭ�bq �+��N4'4yt6��s�Gm�J�d��n�B~�v{w�H��^Kދq�*�tz:І���.D�$�ke;�&	_N�M���ջ%�ke�`crѪ����
)��au�B�/u9��*���,�\���D�Ԗ�����L��jf�G�I�\�7�%�X��B�>�'u�7@���X���x� _�us�c[�N�=�Fm.��Eh��c���������%W�p�㻝g�}\�#5i��-Lz�e�U�X
�eK�UߛX���?�х�'s� �U��e2'	����j�m���R�rn=�H�����q��f�6��O�خ�㍴�V�&�a��Hh8��6���%�@��n�1�kH���M��v$��Y���u��}*_3��˾g㤌��ý�S��*�l�������N��lY��>���Ь)p*V��,��$e-v|��:D�PK�=��E�|̞�;P@�������X�=�!E��R�(������%'�-�"z�EH f{m�M�\% o),{��-G��������.�W������λ1]MЧ	y<F��A��ϭב��R��4���WvK*��)�,E:����056�������7����]�#T�Č8�{@f�z����HQ���#%Ԉ�1՞��U|��9��؃ؠ]pA��
��]=*��krP|U=/�(t�~S��� n13N_"�'94A�a�H �2�1�
B�+��?ӌ�:-R�.f:7_r"\���A6�<���7zKM�OU�B���lO5� 8!S�����Zth��OXIh���H�ǎ��\9RF�P��06LZT#���L��Ͼzh7yœ�<'A�X�*�n@,͹@W�Hڐ{�s��&	��k_C�t�]57�,��"�u����W�4Ҹf��(*7a�h^w���r{�
<��!yD޲��n�X���{�k�����L4�6�}���=Zxٓ3XlxV64EB    7b0f     cd0�:��VT�+星���"�K�P�������4a�������W��Hj�6�4Z�DЕQ��jVz6��ڗ���:6�T�����70�z����C+-�X�z�u�-D���.	���m.���[&]ԒNӲ�xdhy=�P�|���+g	$��<^���@���[M0�C��Y��N��������>�4���,�����Ů#��ҳ@���0�,uם���X^8Q������њ�װ��5tźM�Ǵ4�N���pRC�	�u��.{��)���7T�p</фtv�]T��4��XH�$�?����
��Dw�U�w�Y䚕�$.I��(yy�u�3���k�L�d��W{�Ε�=��"`�J�>)��b��L1�.WH�]����2U`C[��?�pQ~��uU��P�X��ώ��]Q��ZA�4��^��y���x�r�s�
��x�EFs}����^w�S��vis{���o{x���sw������Ǒ|�QlQ�>�ê�L��3�,%˚��	�놟�&}�0�@1Un���m6�=��<���x%B��_��¥sN�^�a�c0��חz	�� P���/tQVs�k����c1�1�c��_M�'a�3�)��U9�	tI�5���W���z�민��H��b'(���) -���=�<z�C g�t>�����x���ۦ�Qx�:����̯���Vt�έ�κ�no�EE�vm��x������ݽq'�Z�>e2^B�@A��셓���M��ܚ^�q�Xd�x�Ó�����*a
?�B�$`%t��z`-}�!�fh`|To��C�d�����k�)L$���ۺ�	�1�J���J�mu�4��7w50�v(�{X��"n� ��(J��]q�
���!�$��<�=�`��h�*�,�A�uf <���GިA�Xn��-z3s��F�o�Ql}Wz�TĚ��3�^���H�!��h���u��o�א�ķZ�U:�	�rC!W�
~�jIm�ك�|#l���R���S���0#������gr�5,�:\M݌��o�R�ǌ/��~[qz�-Ԝ�ͲM��vGnB%���^j�~��f1�!ބ²
��V��x�W���x��j��+�._�-Ui�
�Fbق�0�(���璪^��;��qj�X�x���٧�%��7K�Ɵ.1RN^N(�M`��xG������9_���^���oȫ��0��*{bZ9yU&�C؈Ad�>�؄����m瞴k4uU%{Oٸ����ѽ�p��,�Қ��o�ԁ
�b��:�1����>�Ҳ��ϐ�&1��
�3A�/�)JL���շp"k�H��\z\s��|��[����y-��8�&��sn^�c+%�w����-K(�q��`APYwK:b>e� �V�hl<'rXx}���4r���$J:���T2�=�ķ���;.�R�G�o��k����k��E�B�J�[����zw۩�Y�$t��	[� �MZ�T�D���6.a�y]"l��!��o���D�-����*������ �M��# vf�˳��s���	�;he���D�[/�s�S�t��^g�0F�w��@���9C���, �����\��6�y��Ԟ�f�������-��'}1[K�m��N���3�5%m<�2>��_�CYSc�#���	�LI��A���U���$�rC܆Qf6�ۙ����A�=.?�>�����Bb!�ȯ�em�Q6g�q]�R�
hA�ʜ-�@AD����A;�"��iu,�?�a��)��QF��������i�Y�U����Y��rF'���F!0t/���FѬ&�N��M'��z]\����F o�k��O�LD�[?�4��'����˘�no��ґ!3|t[%�������~�f ���+�Q�ƺ-L�gEԑ�=Zd"6���(�^O�x��������M-2*;�u�e���A�t�)W5�����o���f!��V��~gi!�Z�~����W�X,Q�v0E���}w�
��qI]��d�l�@�]�������f�WxiEs,${��2����+?�xR{�4�%N\�-�*��Am���W��p�!O�&2���� !ͤ
�R5�%6]c����,f��isiT�N���v�&8�dQ�)����ej��4�Fc�����s�����1�;�0�Y������Df$3W{m���F��Fk� �\�޲>�'�8���^�X=�#|��u���\E���X�q�A*��A����L����!~@��7Bkz����'��mȤ}�C±Wh\`��	�����s!;{ǃ��$��9���]�q`�Z�ZG�9�:=�@�,'��Y=b��
��pDG��1:��SX.* �E��<5��0�+?61��J=��S"܁8�i&�%mh"��B��	ƞ7�[���u���l��\�/�~�آ����h��X���~>n�8F.��.��R!��Ʒ��:�ڊ��r���~������
CJ�8=JS9�$Ϟ�ytz��չ�)���ڍ�|7I���y����k:EV�r�ej�@&�.���F����/-���a;L�u��i��L�!�GCr��+���6j%^�#��d��O�M
eb�D�p^ٲ �V���Tb]�}�H�W6yKs��������C �@ޒ�©�g�૬��n F����,D�Υ��ҏȵn]q��տ�R�E=!�Ž�R��?�J��q'�iϥ��i6O>miC5=p#�J%~d�pk^VΨ<�d1'�z�i�Ć��[d����27���
��,$�U~�0��Z��>]wuI��ٱ��?��N9�Y8�7���յL��`��y�O�Y����И��ς��1��Q;<����o&%��i��t�"Θ�8E{��E����k�u'��0�F��T~owJ�u�ɹ���0���61H?ſ�H˷�������m�����_�"�.p�����ኚW�s�0�~��@���S��a"G�Wo�hy�K����A�[���)���$X���`�w�T�����2�� ~�b�lq���wG�=��7���m*UI1�R~���Af[X��m���/gx])�_����W�Z֠N�ot/���ow����w�!/c\��� ���K�n�y�(Mp���Uar�瘌 q�oB��=-��%N|J�͸���Tt0^��R��iCZV��SàY�c�pS��[Cx�^��6)XB�x�HE��i7�uQ/