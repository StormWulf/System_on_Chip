XlxV64EB    29e4     c10�p��Vs����D�)�j�GE�B-;<G�Nb��;�M �Qlas�K�fboR�*	��˱t�"*n���%�,@R��Q���#ו��m2�-�	���	�D=)�������!�=i���ł|��<���s�Ӂ�R�zd|}���;�l��D�R�w����i��=�kHg�w��h�7��B>�i�7c����s���:���H^�k�Q�y���8V�����c��)��9=���~A�w�[Q�N��GSd��n�0>�}������_ˋ�-R�-�N��
����7gܔ�4sY����<��N�Ֆ~�*�A۱�1���	�IB"��@��uj���� J	�7ۿT(keO���&�*��?+��#7ڮ���hsG �VoiF�'�s�2�,a�`�f�"��R�Y�J	\����.���J��Z���0��Tَ��.�.��1=�P�5�ۈB�ֲ�R@ㇴ����N����{6|��j��8V=���ڮ���@Ԑ�ʡEU�|�j�D#`���L���hr�e���#���a�kkL�K<'>G��77�d_�Mp#�S�_�:8!��S��1�Đ�������cG+�����I�$m��)v���#n�?�����(�Pr]w�X}y�.a2z�5ۛ���a��02Bp���>C���c8���^�%#�+��LێB}G	��z�����Ĉ�#��d�;�Y%���\�+o�O_|�_�N<��N�C�=o���8��C:%��M�U�Lk�݈ӏ:�]Dlş�`|́˲Ɔ���j�a��y�.�����{;W�Q�FR\�{W��p-�!�ާ^d���k�hȲd��C�~�=-�s#>�^�;��+�n��|��(��p����t�z����R�SS�p-	�:�a;���Z,��!הd����=���T H��#R�I+�v�AD�;v�:;:�X�)�ֺ��7P����,^�ӯ��ZP�e�Ǆ�ɵBgN))� ������y�|������a�'w�Y^~���ݍ�IUb�1`���&�T�ن�����)��Im�]����"�L�8�{:���z��X.Z��k�M�cg w�V�e�@��x��v6�P4G"Z��	��B��]�_�&�k'LG�S��Z�MZ��!�5l��g��H�-�vZe��v-dA��FbT����mh����[�����V!��/�5v��w��ܞ�p��W�k˗�4��N,��������Ռ�Y�xW"F4��v#*U�\�g�/'v�M#�p�Z�6�]t�I�9���[vX~����A�E>��0Ñ���Z�}��^R!��1Q�A+$�x�'T6��k�H���5U�^4��E�Ro�I6d�#��7��>'Tk�%p��s���*�	SBm���o�㒩9RS��ߙS�J�(��g�/ύ��V(���l
v��h�Fg�}��-��Ϧ�u[� �� 9ƭ���E�+�9r2���j�����Bh���M���K��H���S��@,�߂��1�e��:)��)�M�@֏l�p��6z���PC%m/o�Ox�@~�q�~�-}�|Ƴ#c8V"5ƌ����"�����X��{��e�U[�V� f�[%����94�o�]�0CQ�Q2�_nrb��c�k�O���ً{|.%��|��IK�.],��7��������g)^�y p��f�fJ ��L��{�S<�R&'��V��]z���y�.䶈E�P�#M�����&'Ӈ�!'|"�$�?{F�
f�d���o��ɵ��f��?_~nB�G$F@SJ�b7R��˸S��N�(e}��ݕ(6,��� `0�:�'�@b:e���`
!7�a��'S�Ĕ8c@�[yOpWqYkX"�r��\;wq��&�����*�١�p NgS���O�%���*KB���2K4�	�S�7U"�߼�<�fK2���$�4n+��>r��srA�f�P�2롩��h������H�J���Ɩ*�,'����4�L�d��fyڌ�c�O[�3�S?[ƲE������[Bke�LQYR��p��\�c�&>M�:k���v��o���s����-^��Y��rZ:��<��Y�D� �hX���w��)�2�UG�@�s诠�Gf�s���`�- �����2�O��>��{t#��y���7v����]eo�O��s?$��|��[��q=���zҏ�$�g��+�P�"�W!*.�-�̾�0>F��Kk��	�[����Yet�9ߜ���8��l��K��5��g�b⡁(�8^p�����(���z �k�Co<�f�o���nʑ���SY�����Jc�\�$����=��r��^~($�����'����2�ƭ��q�� �?]���y���|gݵ�E�`�vd0ϗ<5�_��\%�F�7�S�h)�Eq�Y-�D?(}��~���~��k�]ĝ\Ȍŷ�U}���g��d��#U	�pF���A���rB�b�ܒ4ֺ%f�?ܔ:��	^�,�i8�+��wP�З܍�	�j�M[�H��c�ΑL�����P`�ϗz���9-����ע��7�%�jfxPD�|����6�uK�J�K������	u]�2J���A�lR.@bT���q�����Yͤ<�j4�7)��cw���1+X%�nI�������e�(R�
Y�e���"9;�����WQg�,�W5p����z����Im�Y�൙G�C��\�Hj)�дW���&8�Y"[s4���q��Z���}l�?7~�_,�0'jI5{59�/�8���]7d�{S_E%1�����h$�Q��K�g1�}0U#+�6�_@�#����fx��m����
��q��� P�-�餖r6��t���[�{|��)|ۻ�Ĩ�Ǫw�/j�	�>�CV���U�Fr�L����]qY`�bC�8֔R�O^8=+��vzo4���J���y�������������X�ږ%2'�?*�� 1}q�q�y�fO.�7��4��;�����-,�{z
�!�&t���+���#