XlxV64EB    59c9    1410ve
�E�����}���B���H�;Äo���d���d]ԁ�]�,@�R���ɒ�K��[󑓝پhL��G�>���"#���8"?v&y�F����F��(�ߙ��ٶ��f�8g����D�i�\��!|��ܠ����������c� �m(�z��r[�9":r��*�v�����ű�qzv�N��o�pcN�7�hc.2h���Q��-�=�ؙ�Ml�fp��վ�Pren���}&7�<J�d<�0����1�gbXM2�q1=��.A�ߊ���`�����2�753��{������6EB�厹�$y):JZ:[�/a��a�@W�Q�Ԛ�b���|AI
|��s	�P�9��o(w �.j����r^^:�[����Wì����a�ǐ�����W�5��g��hB�=����Q���EP�|i8��j{�Τj�# �*�#��q"����TWe��:E�	�R��$9�{����[r	+�fk�0�:`"���<r�����@R����4�'�eEDc�|�Sva1�5e���J!Q�'E����84E&�]P[{��R�����Y%�s��y���+d�l�"C	c�$N�S� �%��e���#Eݙ�:�'j�m���F���>�;���2dᡦ���g6��!��G����$��u5�����J$�*�j}�Ρ�Y$D�㡲U���=7���E�.�>QTO���2j���cO^o;�m}�>���Gk�-�a$���D<#j�.r��̃�9�x���3W�ӻ�g{S4��*�
ÀV������� ���N�0�g��|�I�W�x��<��
~��5��E�\�8)������ڐ�Oۙ\8zÙA.� ��d2�M���^���!��7���6��..�|�Dx��9E�]�=�1PGs�G�{h�i@���?�q_S:,�A6��k1�O�%U௖�r��2M��(b���r��W�*��X��>η�H(1N�r	�Kl��7�u��(~�f���3��ا�3�v+ �hRs���ZI3r��.l�S�
�9��݋������3x��ʁG"}�~	v@	��@S�,L�4i����`-�.�u���[d�� Ӈ[�}���IxME�y��vᘇ�}p��gzY��hY2�>x.�&We�#�������A�5�s���C�D�G�o*_ėZ%a�����~���a��.�.*!-���}��[G[����g y��A���c��GO���´F�W1|�O�i�U���k�T�ܲ)~�N��+�f�Ъ1��������;Uz���ֽa�N��tM�@����D���N5��Pt�A�Un�LB(��v��Z�'*"����)�&���l���\�L��i0��Π�$��P#��f�s��k�Z5�N���6�c+� �v4�a�pj{���P$���{�K���H�u�
$��������vȬ�;8����,W��1,���%�g�yGY#}O���ʯ�5�g~*�Ѯ��]�s�8l@�L��{�D@d�Xt�%���@���a���,�sn���m�(wU%�-�66 ��O`��w��as��KV���s��Q�S�L���Z���i�q�`iR�i�4���� $���C�H�5[lB�JiG�K�����$���I^ b��1#��H�6�)T��e��]�4�B���*q��(�E�ݼ�(�:F�Z�>J/[�ѓ��
��KH�F�o�2*aK������,���hH�|�ω+�D`[k �
����3$L�⬥��6C��3�ıh<�^�Q�Y�l�����R��s&�'��'F��&h����2��;	�YGp�Je�h���@�p��S4M�w~Q�@���
bP�]�4�Urݔ!�<ƓL�7�7� R��00�I�J~ZD��D��:��K��@�s�$P���ē6�������voOEV�/�aQ�"�b�?\����B����#��Zp�ܺ��,Y��*{+���w��!I(~;��Fi���əf��7K_�s�����E� ����3�}ǒ�r�:�5&��Eu�X�*�{�[����bz#�h���Z?��q�,.�zV���Y3����cSG4o���[G5a��3Z	K;����$7��q,�B��l
�;#r��^w� �?X6���\ȅc`��~�@�(<��$ֻ�h�x�z�W%��=�ߥ�Y�][[���jS!�G��/P�߉�����̓϶��vi �U^
�����-��S�qjF���,�˻�W�	V����2�R�K�2`��W��} g����O]����\�a�t?E�؉�>��߱2^���y��Jz��T��ȦK  �0�GP�&DIle�
/�F*le��1�)=�>^�5G�~�4I����]W>g;4�\�) �&`@��9^l�Q�1\,�آ�.4�B����h�e��ZxD���C�kd��\Mk3�%r>�42�d���4���VG��"Yf�
~�f��eϟ[�H���g!oN�����؂<;�V��i�R,�| o�sRPAҜ���@$�v*��[w�����PY�	��"���H+�d�\ˤa�;<��]H�^L.C��\��x
`������Hb ���l���;/j-����Ç�Fn�S��QE��&R�#����/Q&��k=�r�Om�i4h�j-wܦvh���Yx$
�vs�g��ό�ڡ���Fp�>��ԫ�WNր�����֠z�S?47��rF�-���o�H������P�V��	��
�xf���%���/�<y��!3����h�z("5�_�l|1lX�%��Ey��9Ɉ[��s1&�e|RO� ��T}����W~V������ܰ�h�[{8"��>�:�O��?�^V2���/�������������`���z(j$u�c���<���o�"�2kJO�P!���^S���:�?��iV�)�V�ݭc����xd�2�m4�]K���ӱ=������c�B�YŬ�桻q�{s{�	�=�F��0Z^��a�"�M&m3D�~]-0w��m������}�%'�z%��*����-RN�ɗ�>��Z��B�p��=o���i�6s�~yM���S|hõ�ٯ8�	ZB�p�&�(.��|�g.��$��ւ8�!M� FqB�f��l���wn������Y*ٔ*y���S�ik����l��,"2-�*_�\Á�'m��u�x�&7~��Vq�3��d�)��$�'������H�@�؅q�]���12�8h��d]���+��
��H�C�;�[�s��4I��NN%nl�3�7�^i�R�'T���!�jfL\+�}�q�d`�%=���q�k�ŀ�Q4*�h�u�xeK�D��\<��G|G�ش�Y�С﵂�9�¡�zâ_V�M�%V��(4�Zpհ�3`�h�֗r��d�b�8���a$��&8'��_�?p4Idvv� ��N��0�*�����:��?����" �>�N���[�����2	\�)�����$0��ğ;VU��51�����A3���G��lK"���Gԅ��;f��I��jL�&�;��'����&_���+���į���[��|������=�Q����F,%�=d*�:kV	�? ��}M�bF+mR�y�h��MƯ1���#w閯������^V3�'� 4TV��;h��/�ض�[��ŲfJc�_1|�,�����sᶛ�� ��X�0ŷ�e��s{l�6:�p�OtXdZ<u�ĴB-[ya�x�[���?Ν�B>J�)�Ƿ��l�Z����+�\��
�/�8�hf�w�r�1��w>λ�T��>T��;�?�=���݆�҅��:�M8�Móz~�����i�|���״��~��,��FB����bҺa9��(��Z��!�t�܃\�J�����(ۅᠽہ�P�m-[+L���t�M�N����xWLl'j�Y��� �r�[���		�`�K�6�̫�(57^�Oo9���,�.�Yf���3�#�9���K�Q�:��0���V���̓?F�d�%�� ����\xƖ��H=q?��)����q�M����I�4G%H.�;ɚ%�J\7����P+�g���_(Ρ��R�Ĥ���Q�;���~�J����*�t��p�Q�Ѝʥ���J4�W���%_ߦ�<G�	�L]�������e�.�yX��-(��*i���y�Y�Ց�	�˃�	�q�G0��]�����&�X�%a��u3�q
�+u$��*�u�V�aP\�:���'�c-)��mX6���0/ �7�]���aS1�p�\�։��"�3�`�>fP���P�SYIAL���z�AŹe�?O����
;o��nޖK�_���u�����5���S���O������3I�s�v��n/G~}��'�Z&��9Lf��b�a�1��H8'�����r*W`�J�v���2@�#��8��;ܤ���Q�!ם�g]�V<1���M�ܓx��k0	8�0O��k���-I�����������Nv������e>�n
�T�U0n����o���VdMw=���V���A���ڀ �Tô|����\���K+��
Ek�ŷ� ƀ��R"0=��`�d�KCz�����
8����LVq��v(N��+3�;v�\�k�[ٶ\3�{d�C���C!����v`������bP��������D2����0ט�ja�X��_ގ\�I�:�h�7l��T0������F	����������x冷��������x��y�QL��o��c�?(�P��?���ĶE�Z�~Z��Uc�gPuR�;�5\�������=���-�Y�[��R����ǿ�*����QBM��zS�{"zJ�G*Kj0���KÜ��ei8��iD�Ǉ�~�oM����uf���G�e�����
�ت}�z�pI
���I��Dw�~�f����:7طB��:�З�Y��۪oR\�'�ss�%��r�zV�o��������}i��� �[�8�"���c��B�Υ