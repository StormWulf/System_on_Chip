XlxV64EB    1ea0     a90��I�b��{��S����2�|K2�]D�ni߾�\�7RxzK�����$�R2^!}!ұ,d緄'��	��%D,��,,�V�+ZSy���N��%��חl�g����ۆ��p� ��5mE��%��"�'��"r��"͇����/�B��Y���3XT:p-v��[���v�0y�n��yT*_�6}�/i!��HE/ت��� 0Z\�BCyE�a�.�f�z�t�������w��$0�Q�r
Uc��p�DE>W����{ѿ�b @}E�P/��\ �0��!yS|��b�*%j�%&������'w�ܹ�T�B�;�=G�F���m��6y֡Ep4�f(���6�����s0b��
�-�Au�P�]V#�s��9��h�����k���5�]���G9����J 7+ƓŖ�#�r��;�WC�1v��6�f+I�]ַ�͍Pbo+ Vܜד����Q����1�L���)-�>�{S&�ڑD�L?�������eiՉ���?�����꼈�S���%)��d(�ԓ)�y-z�6I�
�t�� �̦#?p���2�����$��eZ��/Fi��`X2�ϜL���Q�|A3`+�_�ڶ���fÊ�2��@/�y�E���#VKAs5&fE����3N�$=�����fu^�$,� �Ɇ��z���V@�ŗv�F�3W�����X���	zIs�z� [�6H,��;�Iq�5y�	c���)`�]��;vv��q�kׇ���E�Bkw���A�D�e�^�{�1�j�*T�V�+?��о@�K@�q�d�J�r\�+*,��Xi���,�Ӿ��Ц:���Q=M��QF�t��9%���M���X���Uyd�3?o�h��+>�0H���W�0v��E��k,3,6���	ewt�O�Z��I��<�v3D�M����gx�ShHn����	C�.�X(�4�.����f��I6��JZ=� è ��W�Z�tu�Lw��4*�p@��M��Ô%�꫐*�.s��{��θ�����8dI�������a ��" �5n�d�j���uk^����4��Μ�g<�fWf����vw�	������G`�KIl��V�����~Ž����S������mM�3Z�2Teb7|��(�2 ���:N�;��1���w��y� ���2f��3�D�"B�}x5�.L�)����*�*��КZ�?׏͆î�Zg��Ш̯}Og=�}E�l������6�{?���v+}ۺ�����W/����Z�q�Q�~>�@��O�UvM؂�ԁ�7�̙�_}�k��e�{�C��Tef�$������8�����&C��Z����a��81���S�%���Y d��e����4ٟ�l�����C��P`LYObQT�0巻}BG�߃�wC��nF�2�{Ib�r3�H��-A�*�f��sbE
(､���襃�1lM�ugI4� �a��j�>�PY��t)��E�A#/�E��A�,�o/������Debg[�O[���)��F�y��<��tM�:Ѡ�Z�j�K�@g�W:�c����K��{y�&��j�C���)�GN�e0��8Fx��M{pS�Hy�"kj��̪7��yGJk��Q�ob��(b�R�V�m��b8t!]�z��ip�,]Q/�_!^YT�̯��_&��_Ӏ6���7!]���/"�q������ا���_r���aF�!Ϣ��c��_{���I���s��I���\o�=0Z�y,?��]\S�|�/�kH�ǈ$M�~����2<a�RS�zVg�e��]R	�ECh@P����^�E_�6טU�>@�hn`�gp��_���LD���T��{F	�	�z�Q����C��j��t"��Ʒt�����* /Mj0|S�ěP|�=���2�0�f���� ������T�*��D|�2��XB�;�Ґv�f4��c�H �Bբ���1N5˔��.y�+����I)v�S��-3	g�tJ@j���)bXh�`@��K�� �+ܶ[��f��Ǽ��DL�r�7���c�(��������!σv�eAm�@�5�tܨ�E���"-ud����k�k��V���c�%LG����{X�1���p��}Aw���]�j���̊�uo%:x,��6�g.l��}�S���0077�rx����I���t�K��
e�74
��2+�{.��l:q��F��S�h����8�t��>�$e���o�9綈�Af��E���|���{��:�_|T�.�: ��@�F$��jl%���Y��H�y2|�2��Q�y�QZ\��`�Cq�����)�I��69�������'�fE,��r�ĵ'hђ�\:oG��>�~&Z,��No}̱�\���A��������n�@){-���7w0�!�/@�/%c$/����?w3��#�t����+'�PT�`���b�,#VمW�~�*�+�$t����o+�as~~���@������Z���ʳVq�L@Rзq�mi���)�-�ח��ǝ��?�V����kT��X�S(��_��S�
G�3��Ł�g.J?�LH�M���Vϔ�����ʤ�5���1r�sqw��Šv&}��NB�0U���n�bz �`~����Lg��@��n�q���`�8�ʿ2?��hT\c���U�l