XlxV64EB    7a0c    1a20ح�~g���:i�?��R���;�$:u��P��5ykϊr�G��2U�Zϫ~�֣\j�3Qژ���;����Ֆb�) ������t���k5I9�@��!�������) E!$��ALD��wF0���_� ���5��Z��5��%������m�U#�u=IB���%7W!~�{�y�nͽh.�},ښ��Cg��(�&����*<m�G����+Vh��p]x��&�Q��j�
O�xvɧ�Z����3�c��-���M��?P��0;C��=��2q���~����Ei]���A�D	(��E:��Grl?��}�N��^�_�e'X��Ch�>����q/���䎖��HD���!�Kw��>�,��JY5��0֛ƞ�BR�]&ɍ4����!!󕧭25n�|���'#G
�/�h�Q{�L�J~��v�i�0�o���,�U*�U敹���NҰTŦ�Tm��}�>�]u��+��n�yd~(�ym��q��C@f�=�������_p�!�����/#)��>;M�����od[��P��F���r>Q�A&��4O|��\2�rn�j��ڂ�<����La��e�޲9�m�; s���Ƚ;����5;'L�]Sg_�s r�rĪߑu���QuS;G�T>۴BS��D�%;��\1'À�9i�렴
p�@���> i��ղ.X\�)�Z�TyIGUC�8���_:�G�99<����~�Ud�fE��}��;#Z���V���-��x�Js�Y��wm�Ӫ��UV�������|
��&G;��B���r�TU�6��o]�`"��R�Ml�5Zl��-,�����m�C<�H+��8"^ʅ��dYsd��6uK6\x�Ӕ.+�0D�~���y۽9N�.gCx/~��lyu��1���c���2�­,mjh��U���9^�B�/�]&�+E=��Z��6�@	g�y>M�V�s�ެұ9���%�C��X�J�$x��;���,�y�±^
�ǋN{B���ؖ`$��5��3�bB��T	R�0KQ���n����q�N��!w�i��,:�e?��T��O����(�*3���t|5|�?�D�\���n���H����!ⰂB��\�c>���ۃ���y�P����M[$j`E��@�Wk���@�@*�L�,�i.�r,�ʈ��W�4�'"x�N��=���/�����JH�^^"���p�}N���&�u.���{�v	�`1�j��y%"�/0p[�^7m�r�q�сC�Zߤx�F��3�I�����5E�]a��e�"\&9H�8ѻ$�(p&6r������w�]��.6�毴#��!�c����jQ�<���L���b��<Ŝ w�4ɉ�SX��5�v���L�O`kX^����P���,��w:�ԝ_�8D	��d�ܐ��&�"��������x�D�BՃ��}@����g�0��{Xy�/ ��{�����5���= �%�M�7V��zeW�����g�yYE��������g"o�&����]�n�ov}ފ���7\hꊍz`hp��>x�{��=j��D��Jk�G�@%�F� )�.4�+�z	=�gHR%�B��	@����ś<�T>��c� ���aֈ"�,�*M+ ��(u�]-o*�n;�Uڸշ?#�x>��ҲO3�pV�H�L��k�6+;H�aA$G��(���OC�+����N��-��:�uG�X�*��c�nr��9Z]�{\%�E];6 n&>�<7��NJ�d��C�+�S+tM��S�(�$e,.E<�㭄�~�?�-\S��0d�?��rG�~Ɨ��qF�����D�����Yog�)�gפM����#n�(��b��)�fZ����ݺYy�E�������O�sD��M�c�s*p[A��Sҥv�!�k�)T�&���숭���m�dd��|w��ڰ7c��OW�Z�����@�\�
]�+}d֓�2=��������醌#�Lھ�
ݖla�>�0�Uc�2�o*���j��0/�GQ�36`+�*���7lz���$E��\CC��X�I�-�+<~Ws�II��ڈ����c�ŏ{�i�֊��0��ϭB���Rr�c��ȸי��F�kW���^�t��_����ì��"g}���Q�6K��rv�$���P��N�c7(eS?`p�ݡy�
��Vd��M��M�%�ۥ���	���{N�ڤ���\T\���o���eޝ�"  �Ib�%�*	�#G��.��3z�|�mƧ��R��ާ�YH��W�h懤vK6��Y�.]��ú��[�jL`�?�R��9�܎��i�ϟ�R4�`$d���h�oH�k]l�T5�v��T�~?n���[�����:P�n�mg��t�g���֝
^}�W�%M�y<��u��L��9�/G�LWB��i��2k6���� ���4ܒ��U!�C��b���P|��,���Z�pS�V��q1�T��b��J�boo*�����z���R�[:�t�pF��RKSX��=�m�����������"���F��ؒZ��@�E�&(��1�L���w���{��	�M�+ヿ7;��Ö��`6�v*P�f�n1Z������!t 5"��='�r%�m>�.����Du�3F3-��&���b�l ��.c��`T�k���2b�6b��������j���b/�>�-x�p����I��� ����L+��/�t�3�m,�h�1�pV��y�й�&A���A������>��y���)4g��;�����qбj�{K�F0M�Б+�8�>?v5�V�[1�>f�pN?��p�RM&�-�f�b��:�8Ũ8�GFS����
����4����O�<�H��1�G���iTM�Z�{��H~���_����!"+3X����((^���k�� ٥��q���g�WO~���}A��=w��ի��]�佺m"�8�������)/�n�H��KԄ�-��v��N��l�vaΈ{	�Gc�Y��<-�K�^}SFd��ro�|��aS��e£����q�y۴��.�+�r`�BB?B�]�z���Vѧ?��m�4�ȅd�\�4���^�%&z_�c�~��"H�l䭷Q9".�w��*���`�#_�j� sD�{�]�'�ӗ8�+�MG����_�����
�qFU�T��S0	���?4e$�f��"I����{
��w{��Z�kg�
	I&z�q�4�7�G���A��!˶���o���17��!6���o�w�-�}��`U��e�Q1|�W��9�]Tw��fO���{�'y4�wT>����i����M�/���>z����u�oI��eb���4��>&oF�\X��J��nTVE�\g��s~y�էET��GBR��\ |Zb��i>�!��)��0n2�S��zZ5�p���a�y><R�j�	���a���b4u*���QB�z��Ts;B;��S��UKl,��uOK)e�4�_Ӭd{��G���"�'z<�u/πi�Vx9��y��@%(!�e��qc)�W��2ERVO�E���r�P�mڹ|��a�3�U0<�R��<�`��E��bO�o�L~��r�pm[���6��L�!����ߛB��VO0�4�!r�`�>�߹�	��^j��0���3��nw��-4�����ɸ���;m��˭rC]>�SkT�BV���	\�����m�i�~��F� ����]�ǐ�)�.��-��z$�xn�zFx���j���7�j�w{��M���P>�66�W�מ8�_��8�j�t����vLo����S�DL��/��Y�|�+F�L�DX�/���8���?���J`(̭��XB�CŹ�k!J<bz.n/ d'�?�eHml�MZ ��|~��hʐ�����	��%�8 rQ��c>������l�j��2�[�
�����Zk[V��A�_Ǚ28���(;��'D%��ϼ���;8|��D�d���3�i.�~�k�:����P{E �m�b\kK'̤��L�%�i�F��/NB=�<
5l��6�{�݇�=A��L�_���o���~X�MN�T�OfS���� �׊�p)��Ҽ��z����_0ߺ
ᶫ�Sl��/���23���OႻIS`�V� 	=���OВgw���m0|�{�~�Թ<�B�RO�˷��3�^$��^��%B��I����8�Dpܱ�b�B��N��l2e�O�q�G�����9\�?��L�Ӂov86�-\U>��mHc�}p*"@�y�}r�3M<�WT��"�"`'����K+kO� ��إ�ʏ��g����_���W�]gx���B�pC5,z��IR���
�m+���(�*�j4Da�W�ݓR��i>Nn�|�9�0�k��qE �D���ሽD���V�������j#�����Jw�"�޽�3fb��ef�y�}E��88Ƞ~��p��f1�/�^h	�愵bb�4=h�;ݘa[!M�b�1�Kc}��Ga�(,Mj��@A��MP�vb�+V�ߍٰikQ���Q��9�>�.y������N�Ix�T��a#W0��BS�2s'k�Q�m�l\.7yB)!�J��G���g�����v��u�@���UݰK��3_�J�?0Z&�B�n$��%��fcأqK�׎٤3��I���֍�5wN��Pj�$���ռa,��\L�g%e��^������y���h�F^.I%ؒM�*s�?G��єL '��O�wmgoD�X��5[�c̗.�e#��>48\t�O4�T(w,2�~~G��J��������u�c�H�ge��p�O�����~vy%!D&�F 
Ң���;Ed/7T��[6�~>�����`xRK+���<��O�Z���&M�䔈«R����:x2��i)U���"��X̿�%��MSXnZ��ܶ��%�gɯ9�t�����:7b��;�O�6�P�8�~>aj�R���QlJ���\��	ܡ!>g ������.i�-'hm,�*I���M�?Ύ�g>����kl��D'��w K?�MOAT&�ة�'��6��;[��y'w8V��*~����F�
��Mכ�zs���w5�w�8��ݥ�x��D/=h�t�-�%W2V�� �F�!oɜ��%|3����S��j�P*�W��(�g�2�#��N�c����ȇTAVy��#��8bC?	����h�_\�/���n
��g���v�^�ۍ��%-�'{Z��ւs�Y�=�4�h~',mx~f�^�'���Pk5���3��M�6Y�{�_;%��%�7�DW��H��f^�(���x7h_Ï�wi�SlktF��7ŋ��]���b�B���o�{rHSt�$�d�i�j�=�(u\A��ʀo9��+0#�lc6��¾{�G�s���U /����k��9I�z�$�'��>�Q��E�;Q�zRQ�o���R%LY�T۩nWM0��ߗ�"i��YB������5�"B����Ά^�s�3�:�[Q{[]̞9"Y�MDQ?���.��d�J`�����0�D�ϴ1�O��m��
lK���ri!��,U&�lv+���'0B1��m+(��|�xڕ� ��srg�$��ܕC������q)@��p�T��Ƀ�"�#�/��*�z��[�>Gm�qq+�M�#�[�FM��;���u`�(%�?e�A9ٷ&^��=�Hm;���B���IԵ�фF�C��ťb+U�F�o��N�D�K,���CZ�^�#sO[��7�U/�z��ĉ���aj����uV2H�������/.�ω-{-�{�ˀM��y�C5��B�:���dE�UX'R9��}��������J=�(���l�I���9�,&�7�wT>kx懞�H��KL���f'53��ִ|�글8��Vw��ܱ�h!�#lݽ����85~	�����-�akC�FAA���:���k$e:���,� �Dg�u<^CU���y�x$����\�?��}����.&�,��D�MW�&/A��Xne;�Z�Y���=Cz�˳�d
�+�t��=���̌��_��z�E*��+��L�����ntg�a��u�G@ٍ�g%��t�Y�S�W�m32:KӉ�IM�E,�ƌ�ul۲��iI2(���;6��C!�����2a�WТ�y��ޗ��yɦ�G"r��� R�n'X�[���D�
�]D�L18��C��ɥ�z�
�WԤ�]۟�Q
4�Ό�8��-2�R~n�5:�_ d�7��񪁯�U-j_��&m&F]L�pׄ���:(��>p�M�{�TZR�B��N=�"�w��b�ϸ�5���U�
S0�ʑ2��^5PP�L~�fL� l��5������M�B�oTy��DW�Y��f�z_?���u|�5�0���k�K7�e�޽u��l����O��9�7/�H�Bo��{m�;_F����"݃y5-�e{bq�ҢчD��(�@���*�x���qM�A������˷J���9@B���JgK�el2Z(|v����!lY��VH�bW���:U*T�I����k���;M��C��C*&W}�77�n��ޙxv�B���v�$̑��Z\7�$Rz�@��2�	�ׂH�c�<cKE3�]*tl�6�