XlxV64EB    fa00    2fe0������
���7��TB��|r���ܸ��,qǍ��l����w@����d��C�l��R�����((�y�'�~s�;7[�G���2�][n�ID��C'wW{5c�n�ُu�6��Hʙ��=��0r�H�#V쐏��҄�i��M]n��}I#q[׽$����F�$���FtDK�A@���Y�5e:���*������ �����~+�E��cr�aV^I�N��nyu�-��mt�`W�U���c!ZM�����f�/ݼ��A�������k[-ve�KTr8��ӻ}(���T0�oA�%\����Lp~����9����'������/R!��O���xsf��R���:����\���p��o����ܷrz��i�+5}nqw֫��� �\�Y-Mm�=�q�׫Y��?���D։�-=�N[�~��3�k�#�P�������!I�8��06.���p}~�͝�W"���"� ���C���#Na�a:��*b�E���(4�WH�p~�G3���x��g�=ڨF}��ہgg5{���݋�
kխ��GϬa���ƽ��:�B��C0۟�Wj�U�|�jriG^�}Sq\�jh�b�"��b���|%d��0cYF�I�|MX�lHt˩�h��1�U�'�����-V�Σv�f�;�b�*�#����!W�����!���X���`���ĉITcR|�y&����x��o!��o�4�Q�7��/8��͑V�Z�cK����}��'p�r#/m!K�!<m����w�-"0�M,�o�ң�� �~I��w��?�Ҩ�f2(�Q�k��^ǋ?�T��%T���('���O�,>rT�Ƶ;���i�c��N�M��olxXTZ��,��~�Ƶ=����	��K2$K鰊�yҤ�U�:��\߻�J#a^���۟�[��/э<�aR�n���۬_�L�:k���*f8S��i���"<܃�oz��l゘Ԟ#��Q7�i��>�[�}�O���K�æ�H_�a���J]�S��о���_w�S��B.�b�����8�'���Y3^�V��a��yFl�M"Ft\��(��ٓ����|{?�u�ln	[OW��ϕfD�Ȭ�X�!�XY�ti�7�x�v.8�1XEu�dGci�ce�+)�fϋ�S9�i(��!~1'Q읶�s�^�8|,���n��:�z��#�&�����}MT�1�ߑ��E�bO67mb��a�8O&^̜L�(�j3�ؖ(���3��\��-�����)o��E�X�`(�ͪ~|�,ņ͗���Pl�.���@/P�W�g�J�^�S	n�te�Vj�}���x�D�'�w�Ʒ���#p���D<���8k*E� ���2,��re�G���_)yGo�v�k�!���0$V'(m���,E�������+ے8��a���]�<&�r��̖� /�Vъ�K��W�����#ܐ�&��:ض��Asy����_)j����ۏbb%1Ug����;�����{�F�<5�F�i�Q�S�X�\ ș`�i�����k���ʪ�p��.��#�j�"nCB��#�ë��	��z�`��Y,CO� �clc���=y�=� ��e|�% P1��|d�$���O׈����@^�#6y�qŦ\6�5�6�-Q!�ǵ*�WʔN��ZbítS�E���W5��tEs(	`ޅ]�O�nop�I��~x(p.Ϋn��I�����ܞMIK@��d��/w$�V�|���$�3½���1�ĥ	f��#�$�	����@��wʮ�`�OV�?5�^�XV��у�p�;��� ��6�ؓHOr/��fCy���Bs����BsئelZ�k���K}I��_	����XH-^/�%1J/(g������x����A�@f'|�K�8��[Mf΂//,�-�Tڄ�B����z��ܗ�Nf7�b�v�4c,j�Z��=�P���}�*��� �ˢSs"�ǎ���)��/�Q"j��=��`�2��<��pBAA�����ֽ-�B�з�OM_
[rS�OS��袋�s�n�X��Kfؕ�G���r��\Ŗ{�4��/n���~��<Pe���4bǈ<"Ywf�8�ߞ�V��$V�tj��
��ʟ�/8�Je~�$�?.D�n4�>�U����йu�YhO��$��1ʇ,�˲z� ���S��aCxƣX�G�m��:��A����cK�s��"5�=������<L=�+c�s{#p�+Qj,�p<�NF�?ž�cx�]9��@�Jv�>� �K�G�,sR���̄��.KK���~��ad)�~�2�0[7�ҳ͛G5<�A;X�Q#���ˠ�B�b@c�v˾'�1ѯɅ� �k�X�A���D�q�k�Q��K�+�Ŀ�BU�u#�qOw�Z���9��5��7�ԣ7��?2ہ�b2�P5� [Z���M���i������a�L����ʱ���asĈ�/����?p��LcG��*�Z`��"�n|�����ǫ� >Q�.<qi5�/�����)k�U�����,�Y�`��r���3j�}��b���@A� q f�p�]����.�LD/h*��.�2�{�[P���ewt��rN�@�cT=��d%h�4���SΪq�[�����-.򀱨p*��V�n��9��@���[� # �bSq?�����	 ��*y�'&�i�G�vƨ��G���ں�$�O�}�Ә�Q=Uy+���ӛ�5z����`=,м�ҟ�am��ɀ����K��(Q����3�����c��h�c�o��f�Od�Y��k1�jͺw���ⱔ5?+�(�S�0*��L.P��@cm� �Ӂ�rp:d��I�mm-eT��"x_����3�*B��?�?�"�s�u)-W���c|2+�l���!��ub���[��}��;r�ѣU�g�P������z��� ^JR}Bu����&�lC����Y��I�8�c�V����4�A�����ڛ����O���&]�9���f��W�������m����}�T��2S9��*|^��ȫE������VJE[g���Q�q�(qY#;he�uhw>�[�y ���ʡ�.�*!8qa��7�����E�;�	D �(�����O0I�(��ۉ��}�Z2�K���}�2�B���A��H�"ڭ4�����jp>Y3Twn2����*���,C�� �]őH`��UWZ٠��$-Z-e5m̵�e~����j�f2�^�H�Z#}1�<k$0��3U����_x=8'\^�hTZ�Rg��oOfp8�cj��|+�{}qǺ&�=f1��ͣ7���.�v�O����c��Sf>�]*�M���e���ն�-�Hғ@�q�j� t}w�h^= ���V�Љ���Q[�̊���gb���-s݂B�g��L�����|L��8*���ؑ���]|��It%���Xh�_�+���-�5"��v���6� 2�թ��UEmq۬ƛwR"\����?A�@B���eGZaY975���;jn|a���#���[�� H>�I(֌f��4PGÙ��"ɷm�n��|\��Z�@�@��/ֱ��	)�>�eǅ����7�$��޽v5z����Ɉ���&��$��j(���:b8r������͸��s�+uxM����
FQ�EHd�G�n`��p~�[��F{zq�n�u���xc�S����~�g)}'�`�0oxl֑`��b�a�W�0A+��4�GQ��a1�`;���r�D[�N�gH^Y4/�@�@JP�7bD���u��kУ�'0WU�,�w�i[�E�+
 1Hz�*��1ͱ?Ɵ�9�9R�cO:M��G��8�h�	�eOH{_o�Xz�$���J]�� �e�̒^�����F}�c���+V<�h�s�0��5@ �ٌ�A��B�YB2�l +�X1���� �i:q�S����ج���`�De�
�]�R�qh9�^�9K��T��t�0���_3mgz��ޖ>Pq�PW$�6u�,üDp�"����o��}��R�����Rn�.n�n2ۻ���m��('9��}����������z� #�d�������A�mgi�i�cS�j��!?֌6�LH����C�d ��������~�㬬9)��<���Vl<Г �/�ZνSZ�Y�IP�����>�j-��ޭ4���y뻾��=��J���l0�v��0�?!/�MW�ow�F#@bf��4���H�ï�̨"���+�`H._rc�y��Zj���X��-�u#h��	򓖧�09
����c:�E��A��|�s�)"�7F[�6�G�.��z$�zm
9�}dzPz���U5�	τ�����W���X�!
�VK:VC�E��<���}_82Rh�Ql�(�5�XuZ@B�[�3˃1���i��W�PqӤ��z��ɣ���K8Z��ϫ�+Y����0?%iP/���?D��BD���bF��;/wu#��u2���K�.[e7�;l����%v4��]�E�P�2n@�޷)���Yx�i����8��6��5��8�:`얕E�/�����D��Ug�y���������%�y���R������=].���vb8	;��#��0�k��z~�܃�'��!(�n�"t���Dd1"6_L萏��F.�&լ���	$�I%-+ɗ���|ˆM�1�:�<M���@�.$�vR�]��>�XM:���p'���О6��FL�1l��cM��.�h�z���h��ݒ�_t$2y_�t|G������V'�<ǜ��Wj�=ٸг)�".���ʮ����;*��&zJ��/�c�n4�X! �����RG�6$j�|k�S䝘�� �.a�4�t��ǛM|�RrӞ�R5e��nq95Q
I�2����ddE�yWrl��o�_Z���QO��#v���������Ù���hqV.i�p�f�k���kD@W��q����V�'�r2�[���a}�x�R\B�jdHr�E�␹gd�ALޜ���Xi�o�;���dw�V�ʽЁ��)ݽMH
�0>#h����N�]�i���8����;�K<�/Z���'
�����m����l=��,��?�k'�i
�rS�V������[�6�Zf��G]0�P�,�-�Hp>���O� �l�*8x�Fa#w�7�1��!�2�͝�����7�� P�@� �e%�hY�ҫ�[c�7i�J��T
l���zx�c/"F�B�o��A�G������.6��� �;��i�-����;`��pc�r�e��d	�U|5#D���W}KmtGusH�H=�������9���n>��/��$4����X�0��(�趼��'���'CA���%��hU'O�'���U�MҒ��6���	��ή��߇Sl�R8��羝�~~��c͎��Y�M7�e��FT�a�6}�J��L��<gL]Lq+1�%�i#�-�:%bTz��Q���{ǐ1��̬9�3�j�F��N2�Bm��m]�}��7����������}���̿���m�带4���6�
[�3�]2�ڭ����px/iFW%Ȏ�,�u�(���x��:�r�i���c:*š��I�Zo�#�T�
���w�5�_?R�*��+8a�r`��eo���ݬ�h�(9�zRs�k��WW4-��9�/�Wۿ@.Qe�J��� �,�#3�F�iKh̓s-<3~�OP|��0���&l �A��V�)`�W�O=-y9�����u�8j��'_d �/
�G�l:�Ͱ��~/��`�Ն���k��1k��շ��S��� }�m��}Y7��*�"�L6���i;I����m5���]���#�/V2a���Lx���8���l��M��^�zi�B$0P�X�b�]�:�T���^�HC��.�)m��F�bM��>9�GP�������'�_�~^�=q���5r[(��w�u�R���ۯ-�D�Y��I�)1�k;aT���
���rZeҼ�
��xܛ�As��;3v�e��i  �F<yԆ�\~�nT�u3K�P����Y ��_��i:�TuL�:NDfȯFl!q<��H�6��|վf���u��U�4�9�Mx��7�:���#��1�^����ϸJa�X`p(8�x9����Ao��Wp�̩�.֢�M�j��~�L�f�h�M�	)E�G�A��w�1;ze �#���~;5m��Ӹ�,���N��y�*�0Z����RILe�i]�`�@��W�g)�͚��p?�7�&�k��f�~�*���@�'�P�t��Ts��=���@�ks���*7\T��q0�v�z͙�s.�#�|)WaKBG3w;�,��
^����=�ڠ!��Gm����#�>.�\>Y3�"�&ӐF����8�8�^����W�,yL�#���Bշ�dcZ�����S;�G�#�,��E�'O#��l�J�e7ȸ�
��g��)m:���h�ҏ��H˟m �9��l�ih8�_� �)$�$�hʩ�c���	M��:�ֿ��og�}bjh F�f�$����T�8�֒��� �i�Q�K�Ti} б޳E�xI��z{Ե{�5c7��УI�1���݊�V�,��f"�eL��U�O,�ǈ���u����@ٰ�������{��ذ&<����B�TĤ~���س���	ˠ�h���@Y�N�/�E���A[�y�5Γ����
��<�j:��U֨�ꢨnA!��d\	�Y����r�܊pWY����Y��k�o����d��Ŕ����xn_Ф�<�Q]T��vL�����/(љ���e�S!�L�4�dRwu@>�(6��DY�)zaH�Qg��>�®3��Lf�G��VgDk�j�ݡ{|:�[؟���:�jd`8��Qv�<�!3�Ah.�DSn��a�pfv)�4�YI��HB�%��_�KFP?K�֍
��p:z�Ū��-�ܧ�h�a����62�)��#9ZA($N)L�b�PEP�U�,I(ۍe+��T�S"M�����2t�T�ɣ1cmV|\�����./~��M9>��!����Ұ\I�wܨJRs\�vϷW�,}��XC��,�t@鶩��s��]�={����<�ns�ᪿi�N�^�bX��U�$|f��v��g���H���b���Q%���UX����ĥ>��u�P{i�ҳ�P�n��:؇<��88ں�2(�pŴf�V��6��:�G�p���z���V�8g}3G ��}��.;.�v�_���c�	�� �@�nex׬v�ќ�:\��(Ô�3xћ��Dt������t�w�����NL�u�%�!�LΚ��ئ^qQǅ��Q���߉X50z�O;��Oe�GR(vG~F�Ɠ�2S���E˛���H��C(�G#��Na��<[7�n�o��k�V/PCiD̿(0�Y���h��B5 �5]�42Qm�c��i����8~9'��?�eA�4R��Zw��؎e~� ��M�W��f%��v����c%�@�;70�r��\�x���ұ����T&�!���A���N�{�s�I͠)����_/E��H�����4<�?!t6���KKlߏϮ����e�O�H+q�bE��s�������Yyxڽ�_!�3���4�G�64�|s��zX�UT傰\	���rTr��D���>k���T�p�+�z�52�'��Ԕ��f��2�h��s� �.u�r+��@��H��ӉGe�Y�-2�����$��陻d����!d�O1󀗱ֹi��L�8�oŏ�'���Ie��ٹ���̪ᓅA5��![���p]�eW��CH���uέQ<�?���k����	ࠚ��dY[�[N�%Qzfi5n��j<�B��ٰ8�?���A��sQq��:�/�-�aL�/���,:��j~��S[lh��(9�J�)����L<���Q�� 
Ԗ9��8C��1��8������E��:�S�@�̳9;��V��7s�7�S�S���Indܚ)4�vu���u�Hk��I��������Y�D� ���z_!�J�1�����Yqi� �⧈=n�nJ�����o���J�[*#bG],B��Ą�%jߥ�Ώ��~걓EΨV����ZK���m�@��3���6L(����3�O�5�ih-+`�TzY�;�$�|�I}u�����@4��&D�QU�����*���Z53�
�#6�`&�~���c�s��1�0'��Ȇ�s,���YJ�����Gdz�w|�]nE�ߚ·�>tErTc�oT���H�{ #���&-������F�H���|�O#0���:�/-XS�{�}�`e�0Y�����k��0]Lu�w���T4�����F�K�-[BJz��G�6�BF�p���� .	Ezs��u�9h����*�9��m��ҳ؉e0)�!�ZS�4v�ʶ�kQ%���U��ЯT�@i�,	��)����n7A�j������Ο"#n5(�)Y���w|']Y+�U��Y��-��*A���cGJ����۹_G�L��^�����h���슸2��޹�pm�(, �ТM��b(�H��v�8�|pb/%,ީ(Q�� Qv~��}�BA�&>��MhѴ"o�2�4�i�ԙ��8�j�_)-�학7����]�ɉY�cOU`k��R�� )��:Ǥ�OحJCGQ��㓆(/� �MH�����P�`7wC�=��/w��L@�'E�.��=�1V�����#�(�:�nvA�S܅�Q�?Կ�4�I��
�
J��m_H;�tk3e���Ŗu#�٭�a����N�U͠c��J����p��M����(���I&�Vo �����0���?�r��fy�~���k���g��y��>�PN��ɐC��د.uH���v�^;��6����S�qθ�/�2)o��j =�/��a�$�w�?�MdFՅZu܋��I���@�N��/<�s#L�"�S�������^�2�9Ri�R2VAՈ�ݱO�����
�zJnA��9��TS�b�À' �E��c�n]�޳�p���*���� h�?W#$���[&��AZ��B����X>:vO�W�ǅ�z�ˣS���ۺD t�dB���u�k�D@ہ���J?h�MV�}_�;. Kt�Q�
G���Ѥ�8	��e�uy ���q�fR�	�7�ut5f�|L�n����Ġ�xЊfl��i��M�0h�����4s���#���Х@�7�l�`��ĉ�E��ʆm,��B 'B0��V}8{�� �;��SW�^��ͳVt�����Rz���4��#��n�����Jf�L�Y��r����>��F��F�Rj~?Zl]B	��-p�X�w=�S�5���A��0�h��u��{��w@��=���DĘ��S~�;= �����,�\�t,�-�$"�j�'��2o"y�0�$�����o��ة��y���M�c$)tP�>2]S*r;z�� v�Q}d�I���3����z�s�����V]��b��b
��'�YiwW�4	�:Tt~��p!O��a$���(�&���i�I4f;��_�l�ǵ�-nn���L��w7eR�6��"?&6#Nr�M�̠ȇS��T�CY�V�X�3C'Q�J��+��Q͒:٘J�y&�M�︹u�7�����V��ޞ8�f�x��պY�-�4��aV�[U`+c!�?���[O��i2��yXf�G䒓�|p{����!X�a�B3�o�+DM$�.B��-C�x�ԡ�9��+m{��F��5���7�̗� ����?`�����Y�gN�����FK�����y�G���0N�7W!�7U�hp�� �[�<��i��/�;�¾�����׉��D�9�!�5ܼ58G���P����X,����Ͻ�t�Z�YkJ ׊����l�Ti�̥frm1e��N��*f_1&O>��x��4��oN|�]zLf����� B�L�o C���*[R&Q�Z�NB�Pz�c5�<�:N�6_�i�b��ԁ�XS��<��&k�w�$=�/��j��ѩ�d��,�S��k���h�b+��]�FG-��#��RnAe'���H���{����XBO�-J'�	�V�8J�x����J*�b&�Z i`�-A ���x�	C���S�]��8�	�'_�S�p��v�'�Ʊ�ӌB�j�a���ρu�H��\��-�!�ŜKx�i+��8[��!���^)f&�f=,N��u����4��#�0P/됅>�++X1���S�U�J�m���p��^�6�[l]��%DR/�Q��m~�1�Q ���}B�.�F6�����iF�^��h��Ě�R{2uu��&�|q���lkvi~/��͢�:�������)��~��.y	`*�.�-7�[��P'�T)J�"��7XM���	��М	�Dn���*�(]i|rW֪������8�&0`zS9��qkI���w$�O	o��I|r�,��-�g���<���l@�H]�l�`S�����S�ٓ�%�za�=Ё1O,;�d��P\g�?�KkaY4�� f��2D�r�o�&j_��Dޥ��],��4���7�����X��En�Ó��lZ9�/�Km�ܳ����)�gQX�ʦĬ=�N( ��y���S�%yp��
k)j�dSS�X7es��d���_������u��)�q����RMy�}�׊��~��/�Wr��D�u*�<n7K�^�!������]��ODl�|����Y����S���d���%�xi(�!�kP��C+�_lhܮLTR���+Q�ϛ���Ā�@��l
s��O�v8c��kd�xOP�D�*h^z�t���g��<0h=�+c�A�H�4�L��:B�ξ�[�@!��,O�)�"�q��T_�}��;�E�!;�4�&�Q��/�#=�_\K%/�����.Ԕ��i��o�Qt���3G���9�\V����15�+�DTD���e����PMvh��@J5M�� �K7��Xc�:K
X���� ~o�Fo1>H���c)'͛F&��Ro~�*g8���:����s䣓��,ba7r��C�LA1�^�y{)6+Y�k%<ۢK�
�r�!�"pB�o�
ۨ�������GB9I�C|j���u.�@!�Ќ��s�Z	�*7�f�k 3d�	_�nd4���\h�[���(�(������P<�o�=p�2�<K~,	��� ڎbz��5u!`?w�$_�b#n@J�V!�F��y��#�J����Om���v��9�-s�I���M��iS�zu�~g�\���F���W@�R:��0c��{�E+q�O����*�]_g���i��	�8q%���,�Eᐾ�sׯ�A�؉�?:$�I�8*���bv���pC[�}B���*�I���.'��JV΋j(_@��IQ���;%�~���om
�fn�PF�+��A�]�L%XH4��Υ-� M�����ʈ��tn��m�J�+�z��iy�u�E�/0�
�����PʽUT�tW#�Ft�������N�G�FO���v��1��?°��!�T�g�v�\�dI�`c���~��0JBzSVkϔ��G���uC����s�&Q�_��i	�<���u��"�t�s����$��5N�OGڨ�ɳ�ڿi)�!_���'�A\%|�� >��V�(>;�3�
a#1�b�}��uǁ}YV5�9���xj/��
�z�����&=tZm#��]�C�kK��)49��J���X}���%xB�)��0�"�R0���v�
�ZK����f�٥�.�������bx�#�55; �&�ơ�I�5�L�IC���('���0�MҺ�=T���4	���!e����2���b{:���7�Aʗ�l��=�Q`/��sCՋ�JYpޘ�N1��6�0���ӄbJ#Th������T�y��D��j�	�3 ��Xx��z_��<	/e��_��-)�5����ޤ�J��?�I�Oɢ�Ռ�N�q,d���袘@]�u���Y^&y-����(�C���S��4�<�c_�`h1ɦ2f����X1"hP�Gf�$�q�>�B�!��XlxV64EB    7165    1740;D�n��"�����)������~��J|Ɠ�[[�"�Y����2�ۉ�$��T{����`��𮜨�}�0;gy������Τ�:30;%�����#I��5��m�JLc��l�!����������8+��`-��Q.5EA��&��p=���\��pϳ������~z�5ʹ���E:�1Y47����~+O��ݐ����ɒp�����,ڪ����ٞ"w�����\ad7��w0���HX�<�!P�i�G����6�0oh���kZcH�Pk�$���%˕M��8{�ex�+:q�1�L*�$�Nɘ���n�� �/ K��E�upW@����Z�X�.��6��оa7���1���5���	�c�b3e���y�y�P�I��]�wr�⏍{�π�����SR�j�uE�U�k��ޒ�������r��c��
ÿ[��u�+�hȮ��6�m�Z�+y
h�1�y�ߎ׽�X�n���o��o3B�q��S�1f�F�u�Hz�J"Q���.-�ȉ�� ����E�l,�����m��}M���سN����"
E>q�����~+#��_~ x�W�&\E�aE#ɨ��t��=���2�n����
M#1��Y]&ݯRن��Y�bSE{��-e�L�I�7����և��!э�J���~U���
f�Y�.�i��,!S��ƛx��3�����a�����!�if��bQ�)s���+���Ƞ�V������6E�׻[�1[?I�<��pH�a�x���բG6���t�%��A"�'�w+ �j��#�#�7��YdJ`V��޻�Rl��!�>z9.�N��W#!+�LMЅa�	I�V�WV���1P�2^�cv��*Fk�9��u�ֆ�g�_n����,�Ǻ#-?��%6�Q��]���)��=�9U��z[X��cHt�A��80������횺�i>���s�ZW�4k�y ?F�Y'�b�T:�8�@��L�zʏ�0W�6t�a�k?^���ED��~�AlW���ʛW���p��A�ݸ�)�u�b�A�N �oK�>ki>��s�_��jD�<�"Z��U߿���xD���!~<�^tI�����������`��;إA�*Rh�X�������[X䆄H��[�s4�nǦT^�Tq6��&��>�x��MI8�ש����t�bZU c��Ueb -�2�إ|���>K�o{M��#R�3|.�&ěe9�ฏi�D��Z5l�\����N�R'+A"�p��OZ]J"�I�	�.Qu�VUh��Q�<{��%�����j��.W�(82c���T��A�U	�UI����̏�;7g^���������:/����-]���uc�Q&\϶e�y��݋�j���OF�h�8�7���ݴ���F/d]b?(N�����a�/Zg;�lzO��p}%^3?��M�Q��������(�wPо���" �L
z#���bZ�݅�)�W�D�_/��Đ��:߼�U��H��9��j�x�d�N���h)H|HrX�R����.#'�Z���Ř7a�:t�4?*��3�J��C�IM�+89��5�܁�^&TN���&��|��E����Y,��\�+y��@��L�tX�yHl?7�	OU[8`���4��i*4�+�������1|�4+(���f:�em����GN+�F���@7�������!���y?��ڜ��ŘsȄ��(�}�Lu���ʮ!$�0*Y�ÏN���޺`�$9�*��>�Ol�&�1��aɈq)��sއ���jEVS�~��Y%�I�o�$(�J���q��~/3��=#G�`Z<���YFi��9�&K�/��M�}�U���N�pMw2(
�����ibI��X�����Y����<�7$�������8��Շ�:�iR�	��v�^S?4�D]�ܘ9WnRkE�A��7�<�⦴��/����5�CS'�C���1S��C3Z��D���)�MW�Y����K�׸�.����B�2�A�b�x��5}b����}ܚ/v-Y?-,���GC����oW�U]w�D���[��e�x�>�4�ۻ/s�t��=��y�� �ƅuxi4;�I�&,�lvס����_"��\Vn�v=�NXS�g��^9�Q���g���Y$K�����8�c�`��7ez(S��D�A���(������-�h���7�Ĳ�a��r\|f���g'�2�)����Nd���Y�ީ��7�R���?�=GծZ�vT$̬ǫf�X��R��Vb�e+��v2�C�²+�-;��^�B|��6I��*��K�qE:t���N�]~j�W m]����%=~��"�뢋��J�,�`˺{�X�gU�_��
��Oa�w{K�o�Y�!���Z���5��Wb�!�v�[n�<�#y���;�7�F{9�-@�)qYd���Ew�!(�[� ��x[��d�ˏ�N��5-�F��'E��n��¼�a:5����W�Y�3��y�uoE�_	�w��Ŷ���'��7����3�{5�˶x,S��i�kp=�K-��.� ރG�kjU�w���D�6Q�s����{�LFIM���_;��ofgd�PTX�m�7룫@��F��E��ϨNRj�!O��h1�܆$������"zӍ�Vw�Ww��$۝���HA�={�؈����3���8b�woخ�K ��밦���I����T1{+\�2������	u{:te?g�`�N��\��%o(�Õl�����ԅy��]�X�kCIT5w"ח�4��$�� ���.X��{����u�� F�k6���M��a�,�Fŝ�&����ƅϼy}��;�ʮ
���JTU�O���P$�-<�n.^ɐ�}w�{ÝX^>��w�a<�])��T�W8V�u������ȦOu�J�\\���+%�Gb����U��MG��#� A~5���)7��&���� �:U#���.�=ksy��K>��S�����gV�m@#�VɌV'A��Z���Yn6�,R�9�fW������w˘��A\B�{N�`ˏ�o�/+���f<NxW�������d�/h��W�x�.h	��[b���W^kkfI*�p\��\�[x��\)��]���ѡΐ�?� G��,#�g����=�h�[��	��Hjg��׸aAY� ����p��ո�fZ���K��G������֪�]���:N��k���cs�ǌt~�oe�I��0*X�`=�lb�{�1d�({���EO<A5T��F#�S)&���B����v9��_�� "���<	9#���6�����y����\RX�C�}@ W�Rq&�o?x�!��l��'�g��;��B�t�~�,xT,߻rX���z:��V��^-�ĺS��	2/�T+x�#�~�#<�غ���,�~��v��u@����'����^��� -�{dzP%M��KW{�����E�M`E����b��.�b6:oO���+sL��UB�p�l���?! �Y���%�������EL��Z���c�����"��D�S�~=伦��
�p�p4-�`��.N�ԅ�?�i�	�����z3�x(|_!���-!.�٪��ǵ��̋��/K�~�e� )݇Ҿ�������NX��}��;���'�<�e\���[�[� �:Xo�I]�EFg����!b��\إr�g( 6F���ވJ�2�Ȃ��5�{�!]�%��G�/C+H��>�џ�s��v~4=�%vI��m!B5��Ƙ��)��iD(x#&h�$oY1ޅ������v�Hg�%��J��Z��@�&Œ���dI	&
�L���m�^�dC�����ixJ�Iɇ>��c2y9�f�	�|qN5�'Ү�L�\\�o�>��:�Oݜ����2���듬�`�x�K�q���f�&Y��Ȁ�(��M�� �^��@Р�w�c��ou�=�t�J�S���
����3���� �J5n�/v���o����X���N����w�f�r�=1�{#��0���V�)"�u$��dه֣���=���l����5<�����;�?�z���,~叉�@߂��oX�䧙�((I��$� `o��8x'f4p�Ł������^��pR�_�x��h\q��!�5;��<�G
 �&P�P��Q0HD����2M�Q��F��ўR�$0�����8"|X�sYC�b~�_ڵf)��[�(�i#��pl�L�1�_T6���cc_S-�(�}���� 8ҝ�[��h��c���BJ�(OK[��|⺸�9x@��L��\��<X�	i�
��/�dW��+oRt����X�,�R���X����_�C}���j1;�F�����
��Մ �ٔ�?A��o��(K����C�6ByB����$E;.,�v_(
7W|�.�w�c��R:U\���n�|�?��N��>A�ѷ)�yw��x�� �=Ré� �L�;b�(t1h����#s+�����fOx��h��1�:���GEq���]YI������$;�F�i���!�4���Q>!@���Iv�BY{��=� �&wUZ��>�`���I�"#9��W�q��z,R�,*w�s_c�!�&����,�wr�Z6�*�g�G`�?w��d`����}z�f���0I$�@���qP��)���-K�Pl�a��k����"�������^�Fh9��ȼ�g�%��}K�"ĀUQ8bޕ��w\r�aed޲y�a�¬������|�P�ՃxV���r�b	B�h�wʾ�T�v�]�*0�ݢ�_v� �2�ʤy��$��|3=�H5Եfm�/H��1.�?�,��)Oۀ�[s�lD�'cͷ``+�0mH���\��Z��\��\oLI3�9�۷)��Wv��Rʅm�6�(6l�F	VM��a���7}��C|�Tq�myG[�S�'e�  �-�wL\cNq��`�J�%�c(j�����2��8�ߢNWbOy���rW��l�H6�Ǐ�>e��7(a^��p�;�ͮ�@!(�	V���h�Ԟ	�<'u��y|����
Jw*���1HM?-&�40�M?�/r+��z���oEO�bgV��į�� ��-�@#<:�{�V�-�.�Z��I�M|�D@o��""�:W��/t��+��^�Q����#��f
,��]�/�{$����V��h�|������m͸y� 0%|&�d��D��MV����x|��I�l!�����a�]	n���o�m&��E�m_�,J�3�-�"^��84ׄ}���qܗѲ��Ή�h��x��B��U�Ј�wHO��G<�J���q��ծ�A8'nWǖ�� l�<�0Bmh��S[L7אp�n��Υx���͖UM��,B�I�Q�P�(Q.�U
O4�~ݔР+!��藙EЪh�/���Zq�cG��g���8�sDQ���^"�;�\#�(Cܷ(�0�9�Z�?��6^���#4I"�7}.<��KP��%i�^}ȓ`��H�@����R+şYD����VsF�����,4.����ϊ����<'4��C��/$���j10�u��a�����:k�%ﴯ���d�6H�V�Z��ɔ׹փ%V+��z���|�g֫Yq�����Q5<𜽃\�.��i1�(S}��j�Y$��k[�>~h8m$W�vh��/X��N�_�w�"ң�*t#ڨ�R�)�'�F�7Rֵ�B��1����H%�h&�x�Z��������"Z������d��App��c˿ʤ�S� �+��L��'C���,$>ː��!��f��y&�U�0�GHc�l~Nr�[������>3��b=�y����5�k/�F#��^r�[ԉ�]�E�lڸ#�c��