XlxV64EB    1595     840�a�5|�k3�S�����2ga� ��@ah�R"!�O���?֦g�g�*B�+t��a�fl�u�H��>�޼6��E1[�	�Wysm|�T��m�d���E��o��?�f@�%\�������9���ռ)�s�J�$���
�>�L�P����>q��C,5['GAJ�l��O��ؚp>0>>���V��,��]"���=1�h��(����9�3���<�!�߻�F
o�5>e/6��-�47�(nl%�	�z_���"�-�Zk-���r���nk�j�4��`]~.��E�~�M�����5:�P�@x?�Å�;��h�č�`��X��V���l���K��6n��6l=ӌ��T���@gmL1�C�i��͖�:�Ni	������%���w�Ł�|�	�����v��~}�1ȿEAek-���WN��ʑ� (0�^% 1Dn:Z�.�lO�}����[wt��`�|G�
{t�}�Ч�+D��/��,,�GLε�P�!��m���HyKr�Ɏ������g3h��x����W=���;&f� �P}� �E�/�� 3��=R����}0�g�����X�k��B0�%��y���
+�'����ϴ�ٵ�w�� ��M:�� ��	�;��(��"�Rx�/�j̓8����@�`�=�v(�'��ͱń��H�.i<u�s=�谍͞$d����9��k��Ȩ�������G����UaD�Y��=j�-�M2ג�t�* ]�3�y�IJ��q[�p.{� �i1*�_�7-^G=Ң���]>��#��ᮍyHRyK.Z�N�_$\���,��DK����qǮ6ƺy�Z+`+3S7�\m�_�",wQ��d�@���;m�s ���T��MN�D��
�c��2�D؎�1D_��ʉW��EK�6���S�����&��߽��~�`��P7 ���x���h����,�gJ�d�/��P9�2�4\�Yx��^�)utt)�M����mc��=�#�����ႯwP�nR%�fsz`U�E&� n<�HqЬ�B�sl��4���`�֚բj�E�i��ok�+r�/�i4��	�l��$�^���L��mC��v�ݏ�}����f/y�v��i�h� �{/�8��{YK���������~9�c�=�QRЧ}K��A1x�o���y���&Gb�?
8_o�)�z���8��8ԧhz�����g!���K:I��Z~(�^�1�&~���b`aC]��P��[�M� ��@�T���4�d5.���w���O J�oZ��L��}m�r]�u4:��Sb��$�L��p��2�9\�~fe�s�n�\�$ZT�ۇj������2��A�������9V,�.�W�Kۊ�s�X|jY�K��_˪dd�˜EE�N��.���]��Sb �B��v� �X���;���'�����򧧈����(-	R��M�j�����2~�BM5������ Q���DȀ$b�J�	��5��-Hv(�b.;�� �D��jXy�h�C��Ʌ�v�\�W�� ]׫f6����Wp���1K�@h�BD2JVK� �ӽ�3J��p��AiHK0���P�X����î���0}Zj� ��r@��� 5~ht[
���r�]5�̆x# SA�Иe̛cKyLf�
�(a����m1u����N3�Mx	����'`�m�9��$)��ʁi0ѷ���R�v��lj2���J`��K���DL��3����v��w��S��d�x�轫�'<�P;:1xh'J�ۂ.p>w������:s�_�� �3�J1�K�*�o!|eE�̼	0"eM� 3�\���q+�.}d����7a�!�鐿@NO�M	����ˀ��/�E�6Џ�}�M����nf~�Yr�֧�&����1�˶�?Lqv�L��3��6��&[�eh!Yu`G;�iIy�o�q2��py���a�<F x�>��Pׁ)�uZ���;+Q���w�ƅhT����'Q}/�~�����+��U}E�����q�+��f]�+nn*��}�	��=z�?��Eσ0�T�N���ʆ�������Q