XlxV64EB    291e     bf0]�^���66Z��2��\�[t�^C�\U|�,<�̶5@I���8����z���+(K����/l��#�o�'-���n�P��ƨ&>eq��:��d��R5�uUhGG�)%Ȍ���X��g��z��VT�'�v�	�2x5��j��'��Z�c̏ �Zx���0{�V������_؏��ּ��4$�c�J�0���(���H[�Ԭ7�®q�Z[����#��u���29P�a��i�4}V!���&���ة<�J_/���9�&�j)�X�����!+ɷ/c��s�@=��X�J�����Y*�ؤLjB�k,�7�cȀ���sgoY��J:5A .]N�Ѧ�c���7�̿K�}ʦdM��S}?C�&Ƃ��1?>`�#�p'�)�ىO����iW+����0�-s7��óWB��?���^�s�{��C*r��j9���ۀqvGT�H4�q�bA�+�^��~��	9~
�'Ĳ:C�����
N\��4�i�d!k���T�'�� ÁF���(aHɀq�>�C�����zI�ꉒ1 ��vd?�+(̔'Ȫ�	*)	��U�����ai��Ь��U*�G�(��y䰮4�C0y�aDe5�d�,���^j�}��ϜV�/C��"��7�X��,ꯖ;�hKc5���wј��'���Ĺ8���@�#�H��*ُ������I��Ҹ"mu���^J��/+�<N��ǿ�����FX�֔����+��\��V�MS?��B�&ԁ����<h��㇋��Ƕ���q�(�<cio6��[�uF.�E�L����ĺ!UR%��I�e�ܻOL����A���(T]�������lQ
�6��3�Aj�^V��A�O��Q�yV���Q�ɹ7V5fD�����0��)�#���ac��Z3�xE�=����&�hF��K �c��>����T�1vZ�ml'��\�S��'3]�0��T������\�o2��s~�7F֏w}�l�ة��P�|�x�����A&4*R���M-����~	�%=ӈp�ˍ�7�+[�v�����(��$c�jݏk�5`�&�Y�2�E���.�����$�V�+\�$+���C�h;�d|v�U�ڶ�BNTsәQ�5�?x[�s��"�5������!�߼���V����\s:�0=8f|��i]��q�d�/{�BR��dDO�+򬋤�����54���X��E��Z%��Rz�/K��쟟�!�T�)_E�>�59���R�.�.&k�,��$��g�ʹZ�����N�	U@�i-Qg�ë}�E����գ�S�⌃1��w�{z$�?�޺�Rx��D���u��F�����kr[r�ڷÓ�C���`��M�]�2�m��n��$s]�u��"�_JN��l�]�?���bڲM�P�ׇS�7�x�|a����o��(E��Y�$_{������#��?��k��aU�z��^�S@�&j�F�"Y��Kr���6G�,+�3��B�aEܚ���Q{��#�!I�!l��<).�m�1�(�?ȳ������k���$����BWdL ����<QoƦ������Γ���&]�@ .�vz��B�8C�!U{em��Қ��JY|�;�$�R�� �j0��� �խ��"�rk��葥_��<>��J�i���r� Ҋ��|����v�4����R�.����o�gcR;;���M�<q0���aE�J)�-�ޫx��^+��༈UG��b0��p,NB.�X���2��}�-Z����+��?���~E"TP.��h���;�cGkiJ�n�m�JE�+Tg*�º�k�S�X&ؓjT�-r�Ǔ�:r'�*��_�)�Kb��gJ3�������;N�����|veO-_��L�e�(ӵ�N���+`~�Z�6�&��s��e3]nD�(��^�wG=z+�X��:o(�g����Ii*�����Y�%�'c����>$Wf�oC�����O�6�ǪQ���P���jIJؼh�b�>K�g���K��X�Yrx����\�D�+��?���E�p�e?�ȵ�&�u��Ȩn	࿊�Aǣ`�9G�1������\k6�̐�@1��Cڅ'\�;�b�TO�ć�'`������ i/,$�f���[�����+��}v�?�e�8�����T=&��)����h9^^{	F�~#ZY��E7\8�g��!�]ЉPk&�q~����p�"=*Ȓ�.>�#����5��a�yH��c�=��C���>��MH��y���J�X���X���F���TĮ����.�t�OR?\R��#�u�B`��̿������G�o7������JH�i��dR&<^��:�^���f�/E�h����*�.��YLGuk"QVm���C��#fK$t@4Tr�| ugj$�}�c�ZH~���s*6��R�s��㠘Ȓ��j��Y����?�S�ƿ��;@�q�n?#��O]�s<p�(�s�!Pt����bήH�s�2��ɏh��m殾^�.e��M���1�����̹�i�O�������L��Y���e	�?��Z��Eu���]�0ͳ��\J� $`F����HVlvˇn�A�\Ր�t�A�M��m� � �� �%�	O%6i��
G�ê>�]�MeD���s8o��6���87����y��,B��ů�7f��Y?3�J�=�ٴ����[���-����"��© 5]�C��De����4+��m<>lU�7 ��`(��Bܠ���|���L9�����4�Y�0r���&�F �-K�N^�@RԐg�,��k�������?ȃ���`�4����XY	f�gnxJ��Ɯ�w�m�.���-�a
�#�+�g�i��7ʅ&UxFh9�v� �^IV�TY(�<O��<�`��T�t�2J궍�4��Ȋ����v���HD����*X���2�-�J}�y,����f��nפa�)�r�w���2��`ν �a�Jt�I�K'�<@����N9J�.��i֕o��