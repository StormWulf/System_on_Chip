XlxV64EB    4a09    10f0�^������S�,�x%��h:�(<�O��>�c�1��;tU��{��=�ҷ�@�#w�T���*A�%��3��AE7SQEe�b�,VG�$U�v6��z����r>�д~��Y벳[՟z�4�D4f�]E��	���P��(��?&-�e���_*��@��@����ǎ����X��\�^��ϗ�&cF��թ�s�2gqjR"�0^�-���)3�����m���3�bi��;�J���h�ꡐ7��*�����!(�@\�}���2�H�>�21[�>[����G�p�D��d^��/�������&�����E彖G̊yuHp��,B�������X�Z������7�,ND	�6������	P��8)R���8WK�@����cT9@q�u�?2�R�^�_�$IC^�xu��awP:�k+�������6��M��2�dq�����Z�O��Mf(�Wq4�n�;�5?/�t9�'��T���[̃QJp�i"���~����v��0G�
�,�˭g �aҋ�:+᧻1��X��S��w:�:�!leL�dx��/e���\���CBM8I�N!�rWT���֖(�9��}�mP�U^"��^>\8f�n�|�c$<���� �>t�i�E5���	�gQ�3�l�d2#x1���Y�V@Z� �(���P����o��X�'rR��He�'����q�H�Z#����
�x������Q�n�^^��1;�S`L�m
]�=�t�Dc?�)���\��f��p*��Ic�&`͋���D`~�Fc���Ȗ�Ə�c5�3oPKUr��.��n
b���7�,��l��u�Ta�΢g���gDC?2��z]:���[%� �۷Ti%R�o���.�Ds�c���)u{���n�&,M�wn����փ����b+䬹Qd����f��0�kz$;� �G��X3^�-�OFC�cw�W�"�`�̼̏��VlQ���	T��@"c�2�UU[O5��ۗߘk�+���Q��2_^P�C]A��^���ʑE��W[���� z����`a�70F��[�h���S��������s"h��A[C�J��=j׮4�ǂW�m�&�䜎�6�;�o��&��!��h~�j����q�M��v�c�&}v���� i���v�K�L=j�("Cޣp+�;�'L.���[\�I�~2D֕U�:;���r~���`�ғ��w/�׀�M�ٳ�i.q��}����S���g�⵨jK�L*�XծR����/b���Y��E?t����-���?��=��I{�v8�AW��П*U6�+�F!��Z��m
(old ��'�Rܑ78����c�p<����=�u`_t���P��m]9�Jm��N�,���ˌ;?%a���4 a���q��u��ݕQ���L3gوh(���U�!��_��%�����?��@o: i��y���f>j֬9�cH��E���dq�S�"8h�I�˕���H�Q��65�vzS��0X��+0�ɿ!�􆒹I@0O,��n}:�L�UH&GO����
�u'nE-��C�S��чy��;1b-3��%�^��$�7S���}��;Y\��������cw���̈́�$���D�*�Y`8�f�y�=7���M����λ�Hi/��Y��1���j~	Q+�/K/�SW��ZL��5v�7G�nf?��G#��q�g*��"��}�D�-2*$$���eq��Y6C
�T��؝��v�'k�_ّk�Ï��h��Z2j7��8�_g�%*�[�88H,�_+A���Ö/��$Uj �)3�f��63�q?j�Ew��&&�)�m��N�,��o�m�\*��!QezQ��l�F�F�S���8d���6(wKU�f��J�z�;��aB�2تs5������@.j��l���~r��WO��oA��n�[�Í���v�$bQ����9�Ξ#;@n��|�{'y�C����8s�dLrp�6�nׁ�|��0���5�(!m��T9ܡM�,B���n���E���=�a������jN`����缨�$z�^�j��)���%Nov��e�c��Sps'>?<�S��A��,�3R]��	�5��5���j�9�r�i� 1�02u�M�L�ڳ̩�e�����Uc!�nȵͱVqB�ԓ�BU�:<t��R1g�]�`~�ᆺ�8����܆vn̪�SK�`�\����7�Sko�v�0j�w~�\����^��Z|Brol�����V��W�� eG�=�,�� �7�#��ĮN�O�J�����rb
�����)�D��L����:��&�fX$�hJ��wf�o�ɇ(����|@�2�z�����˶"�G�s-�-8��!ެ�����YW�����l)H�/�q�jy~��*�����0A&n�
�g}� �\O@hNo�H�V,Iz����W�τ)��mD�`ġ��s��J�lDt�?ki&�."�f�'�?Ub�o<��I��[�p��
��W�l�� UKk�E�7�m���j�d�T �7J���6�]�N��+��R;�x/�H�r���M���N��P�j���_I�׌�S�'������i�R1��c���d�:EP�+�����+�������]Rb��m�anRUc�;�э����}<v��m㮐������a���<蛪ŀ�˓������E:���E�G��=ܰF@�/:yX�7_o�,��c��!g4�$F.����c���g���&rL���j���_���q9����X����6��T1�7��/44�¼����o�ޑ�~�v/ݼ>"'�PQ�,��2U�~����r��䔈#��Kf
�k�a�h��}�2!�Ɖ���.4\Tӥ�xa]:�ґ�M=O��_ю\s�HB�9���ڴ歺�ˆvK�AU��E��AB��X3Z(�=j���HJ�
x'���K��u�O3�����4�n4ƥr��3����S&���� /���+���$vl�;0���K�d��_d}M��o�.j�����}�5�Q�����<������죶��Rf�~�@�0>^OJ��ʳ�����4���V?������cz�
5�fBR^@��LF�Ȧ!)2�c��.[�d����fY�y������'80�-`�9�����Au���	���ZaS�5�ܒ�[Rj>u��e�s���+S"��;c�}����P���]	��8���B%�����b��a@�7z��s�`�$�5�����V��\�^m�o�<�n�/��l��ai� �.��S�K:�ŏ��}�'��ŏMB�S���{n1u�K{�1'S�>u�0�ԍ�5�a��G9�̲I�)-1R����ӡ��xf���7��,��YM���%��:��0�w���=~���q10\���9�?-rty���1Y[��uk�q\ћP�s�$�L�Nݺ�ₛ����ҝ�U���n�o����Š? \�3���� �mMI.�c=�,&ζ��6�Qº.Ӟuy�䚳n�\��l%��x�4�'���,��mQx�`4���<x��Wz�w-.�0����o�y�5[?�F�ً�橭�C8�>��\Ѓ���-�Wdm�7��lј_�����m�? �2h-�̖��3g�5b�;����q�Չ��v�&��������S���<�\��>�������Ӧ�w$| ���3����#@%�s0A�I �|*�
3N5��Z?W����"��Rr �74 �\�.������)����#l �nV�F�L���q-؁/p���,5��^�@Kk[�4��+cUZVU�'J\������/}�p!���E����Ϻ������-Rx��K�൤'p���x��0_�C��ND��C���ww�L@É字�����N�d���7Vf5 ��=����/#j������Bg���a��)vf��Ќ�Q����F�:	��l$y� ���ȧ�>��S3Kb"��5_��^@h�xu 8��~����^�GsR������2iO�՗���Q�-�A�����M�`E��K�:X9���V��]���P�x���ICd(9m6 uA�C<���C~����/9�Y|��ʢ�� ���Dܱ��I��df��h�𓸐��N���3��U��"�y�7���v��|�T`ˬ ���K�m��'�;���ScG�,���=�x����B�"�������iW������5����F�/���U�Uk��:�9�F�\��~Ѣ]�0���G���?�Pv{�X{q��nx��ܓO
a��]