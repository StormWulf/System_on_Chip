XlxV64EB    23e1     b50�����REԿT�=�')��y*FMdٝ�@�I�+-�gF��>�*}��ew���\�X�v���uF�¤�*�Ow�QdT#����ro3�n��|�Ve�U���Ec��u��������&G�I��B�w�%m�֍�;1G-��D��~d��}*|F���?]D;��l��+�ڟ����Lh��! ˫����X�!P%4X7O%�~S���E���Ls���?�c��h�*�=�7���Qj�!Mխ��#�P`��9�	�/b����&9�e�n�?\��_w2e�%8[�*m'�y8�aͫ��B*͙�U��:9���q�Q�<|���	�E|�<@5
�t�������}�g֕3o#�xYa4v�K��g�bܦ($s�	Q�6��o�L�$5@l����DWKmb��޻��Kj�H������'�}��f��D�>��ˍ����ܱ�c�1�7��.w�_@I�9�ǣv��c�P�h{�zn*�[�g--I�C�%z���"Df��zӕZ� �gf~,9�ɣ~��g�;�~w�W�Ox%�Z��,NG@��N��᧚�KR"L?'�J�oO �и#�M�u�6`�#�e}���(��=b�F�͞>Y�@�y��;�h�R�h��kh�O�_׼Ut�g�W��%�B^(r�y��>�;��ݔÏ���m���ÝL��y>�KQni>L$���ĕ����-�
90W;Pp��C�xXY��\��K�R�:��e�����ۙ�N���e����p�ڞGu��}��)���eEձ��Ϙ��뻂|�C��n�X����UŇ�j�vr'��gT����dx���h����â��OǦ� �>��ѩ6WWG���EI(���١�C+�s�;�����*�Aޔ��g,|QH�)WtG�?2\�<�f��O��z����*x�db�&�mlBD�N�ΟQ�����#��Q�e�@OQ�ӎ�?CD@�o���u�*� wE���<ˈg�	��M�}Dp6�h�C��OD���Z���^��3��>?<�T�Bg?٭�ms�E��q���mV0h{�`o�M�+e�A����F�8&��K�R����U��W��/$F!3e���\����,����|�V�Q�!ʹ��@4��1�0x(�݆4ܧ��RUSc��Rk֎	�;�|ߑ��}�"�G�¶\S�@J��cL���i:D���hҩ���z:�o5�<��x͆�������k��)-�c�e�y�˳�lp.ֺ��Y3�ZD#{m��i*��~^���o�γGЖ�x@u5A��i4���&� ����q�o5ᢽ[�Ax�c�� b�����^�N`⟫^He���.*�	l�Y�����_Jb�0X�&jGt��g$�ޝjr1c�_`�~٫ff����c�eO4efŒ�hk�]�Q氋l��O������Nt.���S���3!�bh��aӨA����L���;�ږo-ث�P��k]_�m0DC�Y9���<�4YH�����jDU|�:�=D���+�'���J�p�lK�uڨ_zAn��S �V�%o��v��`CK΅��u�s��H�֐d*�c%=o[a��ހ�- P���B��I��#�@<'G2�}ũ�V)������a����`X�^G�%7hV�fbA G}g˒���R�(m��=O󧍵���w�(���r~h��,F��J^8Ρ����i���e�ke�:l
�P/��!|�:	A�f�u��Bu��)`����%��s�4���>a��,���cs�u����پ��(����#�"S'Ƶ��D>L ��W-M]&sA��kr�c�� �]�z���M�I9���ya#�+j�.��#$�d���?Z���`;���S�`�wY��IG���7C
.����ҕBg���7�˷�����r��y�9�"0 � ��ÂآqF��,�҉���2�l���0�B�h�m�IJ��ۧ -I>y��#�"!�Jڳ�XO���L��-��X� QŘ�Ч���S��~H:�l[D�IЊ�w&�+4S�2�g��������^s��\?��ᷲ��.M;<;�!����5$�	�Dwe,a��)���y��#'���xa�(�`rd��Sé9+�`Sp��,��x���5Kr�l굳zI9GO�+,�}$(��-�Z��w�錧d�q�vJZ�H1ʘ{���e7����&�L����֩����������-:a��x8s�	�gֵx3��3xvZ�����$�N�������D��Z���?�p$���}?s���AZ�.���-
������bx�T�-��Q�#�Q�$��t�k��6�*:;`��q�k=���26���V�O�=7�)0@����o��(#��/���4f5��������h+���{�n��A@	�)4l�1n(��V���ya��l�m? �[�+li�1�D�A�fc�5�������5����S���p��h�!�o�����I��(v�͆6�Ns��T8!G�&(��	�o��o7� B���f8��3'���](`�֣@\�P�� N�r0�(���ֈ�v�Nc�������(����;{e��4����P��,�'jlF�xݩ���b�@��!c�iB�6���'��v����G(1)���G�#�R+�pf�a������=��*y�+~�՗BIǷHW�L1�fv�'&a_������0�i	N6ƃ���[��˨s� �q�F����v�|v>4�X�� �7��8Q+�2�y�G����>��V�I ��d4���T�ؕ�P��Y�q�NJSj��=�,���ԡ���*cխ��U�oJ���%J����l�B�Jr