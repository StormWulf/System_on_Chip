XlxV64EB    181b     980��/�4�&�|�ы��l�տ�D�}�yz��,k''~#�qѣ��tЗ*��������iM}X,��䝲�����Q�
��?x[Ƶd!��̠�+���ee>�h�F��j�s��Z�Ig� 2������	p�X���:��o�-'��#,�LApU}Q��=m�[}b#�R�P�2�̓��HK4m��dY������X�.��'�Ͼ.z4�Qٙ�$����Gf�5�6�hL<��rt{��r��t#��@!�cLg4��EK�`[ EB�c��܋�^�^Xղ ���j
�E���;�lM��T��f#�8vvIѼ����8J��e�-
�B�?�t�F֔�D���4�7_���S9ٜ}4ݩ����FgP���������jC���~Z�a^��~�����%Av���ώA�`��6l���n�<��J�,q�bS_�
u�{F@A ���D�zR������u܁�)XIW�J0������p�s��4ぅ��L�L�-'UB�9<�+K�0�$��^Oqތ���k`C�U�Ù�O�������I�>�>T�|�n����̊��mj�W�v"�Oz�pE훇�m���DM��Ѩ�k�h�f��41Y�,ճB(���cNC�bsɢ�=y���GS�v�4��,o�����Q@��6��F�-�%�H�mk��<˦ag��tE�0���xj���K7m� �WýI5d���uFޥP��L�c~��mvmlb7�n�r��_x��4�i�p��vEY�T2����S8���x�v�#C����,�����?9O,�yJ���A*C�&t�9��O擂-au��Ж���#��H�'���o����P*e[������QT�Z���"�)�W���@3~�E��3��d�����_���6>�to�Sm�	��`�ϨF��h|"��XiSe���qx�ń�B��:��� WgZ�Vft��E~:3�ߋ7���B*A�-�i4���X��K#1�E+��,I\򝩽�Lcz���W�/�ˑ=�0ڻ��rO_������;�g��\s��a"��أ��TyEr-LUm&�:�9�쨋�����v���
��,�08|�by�C����_=I#����]W��� 3/��i�a��(�7L��a�Ǜ|��T�4Pt��y��o\I·1���))��_�?ɧ"[E���p��p�|�V�J���������G���|����šI��1��5Q/�q$,IW}t�y��v��69m�P�"����$α&�l-O�6�A��OLt���!�N�6���r�;W��=G��S'2�#� w/C�0S�Ɛ�,=��/�3��h&b
���@8+Fq^�
<��P	�n����"@���!�ׯ����\�� S�@����?H�:�h�6��F��e|4��������'�]�t��!���Pg�ij��� <e��n��HyY#s�{@�����"����C�,���Ѩ[��5�M��M��N�+�d��V]����.Bt�Po��N�Z��3�>��
j��ap��$l�.*������҄��u�%��,��,Z���N�p�~�Ŝ
N��G��F I]̊s�s�ƺX��_��4�ݒ�ˍטx�ڃrl����K&ʞ�Xs�^�Q��Y��Y�q����8�A~{�s���n3|���>gʹ��K`3�t�Yr�X��N�L^M�%�����p�.���Y�==��&�\$�o�̭��R5�2��ȓ��T�/:��[�����-�8��AR�?
��=�i�ef-ׁ���t�֭i�g3�A1�M!L=F�3M�	�:S	���{����c��V51|�Ö́P�=����M����o�P�+�K�p�bLr*���<)
jČ3�#$�t�"~�f}���cT�J����Sy�#�}���~���P�D��o8��G�WK�t�i�k�q�?u���eJ"�Wxu������-�6²Ț�h3��(j6Q��K���$3�	m�\�00��Uu\hU� zi�V���o0�3}��PԨ��duM�q���F���R��N�d� �y�Qz��%0z/Xt/ �a��O}�H��~���(g�
�{В�;�]�e�B>y<�N����v� ����q����aY�$Ɩ���)�f���VR���H
˵�W��z��E$���	��%ݾ�� �Qܴy���C����)�L����f�>�5l�q��q�M��6����o����|Ʋ�x�iE���4i|x�`�����9n{<+���(m��w��,s����L��������O۫��U�W�gU��gA��;9(����(xt��1���%���?`��r([����D�jGo�e�I1��g~�$_����l���$P�����&�$H�YK���8ځ^�3}��0 �v��0