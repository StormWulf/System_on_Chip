XlxV64EB    19b0     9b0����n��ka�� �� =����h<[���B{>�G�z�)��c���q�[��mt��Rk�d��SbBqzڹZ����[t��1�g_JAC�����r������´j0sm��c�`Mȵ�y;##�:'��\%Ew��Fg�J�/��3�g���K������p�>.�[�To�t�@?�H6���u�`�נ�����$�C�Jd�"e�N}���G�hJ3�1$l��C���(�$���^~J��O@' �d�Xj3\���� t�W�^5.��䐗�$�������zma����u���gs�̟u�T��"�cg!&�$�F�G�B�
�$Ԝ>� ���Pn�d�-,��������zFF�VۆQT��m��*�S�<]-�3�t�tС���� w��� �j�����t�o�{�z�C��o��F���2��L%[���N*ߍF��lLP�aWQ  �V�M�ؙ�V+{�<d�nu�L��4Q?�絴�N��������X��3���p��p�W��Eu�*D�������V��,c+�&Q�P��������8- �IP�S�.�  ����Nq��5^*՚��I��6dp��%���N?=�2�ʃ�A�G@�ε��ΰ���Z+]*@���
G��w*��L>�8/�[P@��r	y�h�v�P���j=BF���i��u�/��L�~3!c{X����y������5@3fȰ��x����R�v��o]��]���;ZZ?5=�T<cm�7~<5ۃȜ�W�e�pt�~����+�kL�ƻ�e�W��O�Ž\��P�Z��8�}i/��M!�8�I�wsw�9>� |���D�T>�w���T(Y�7��y�ȵ����4\���j����nI��V�� ��]s�}�P<�1� xp�o
�+�p�ߚ�k_���Zߘ�8=�C]rQ���:d��5i����`�'3�;��/���4���!���V�>u_M�e�Yv��2׮7�J������!�RJM��n���:ș:I����0�hu0�L&N�ֱ;���j��ဳ'�7�w��5ݲX��6����/�Ƥ���ө��KJQ;�]B�� �J���`I�|�f;��]�Q�hK�'�u��uZ.tfTE��m�v6�HX)W_YjM �z�@A�>K����<�@�Xv�]�0.%��|E����j�qXiI��ŭ#d)IP:xS���ڛ��Kेߕ�K^�s�6.N "^�G�S� d��W	X-��fH�i�a�<�p6�ǷE���{������-��[xR��^O���v��9��D��ܜB� ��y�N>,v��N-�9M7/�R�t�M�AS_�cl8w�e�7w�&dUJQ�F�3���7/�~p[�e��C���p�U
������u�;O�Pp����H��Lz�ܡ�"�k�k�I"'
�e�ٜ���%7�����C/��k|&�l�]��7'
䦴����ld^��\�p�e��r�� �Dw-���%L��Y%Ф��H��cKm�	�"b�R c�;��>Eǃ��g��	}���`Z6�Q�:����#��|�ݍ�v���S�>�ʢ�����@k�r�XB���/#r��`�3(R���?_5���}N7bĭ�<y�i������i 3*R��u�<�`�t���9��d��@l.�����Y�,�b~q����m��[V2������*K����5��{�<�,7����p�@��f�/��Eȃ�jҋ�$q)��q��D6���^eP�)X��l�I��B�@W��މ	Ǆ-��^���Hb���x��������)���	���C<�^�-�1'��K�A�X�M]��/�32�+���EQ��)��;��P���sģ����Pov��R��F��KVd�"�*���@_�uH(8�+I�MO�vT�-�ꛂ^��fv/0�%��<Gc��D �`T貿�[i��W2�v&i�����K��-m[�'���Y�v��f� g?�7Q-F�RY0(�SG���}�_��+�[�Z�̵�L��ݩ�	�l�����)	.9��q��d��04�H��Q�#���Ŋ�7k��L�b8�E��}�A�^��q��*�H�إT`�	{2��O�<9�&H�t,�[�����������̠�f7OC5���o�F����p����}V�J�{ ��G�~×��{��ȯ>Ma<8�!�Lk߿�3v�|a���Y_F�����t�H�&Y�s�� W4�\qǆe��Tj
F��\.?w��|��Iao�N
�*+w4v�M�}/�F|�0O���u��;���6{� ���K��ތ���Gl�ql�J�APs@^�KqG�5ɲ��V' 5�#�"�wq`a��V� �\��[��JY����^����J�����|ؖ�	����JG��rE>�W��b:��_�"���U�x��h�"�y���
p!�`�S�2M���-