XlxV64EB    2279     b00�=�9��ʉܣ�J\f6�btUKQ�瑀M
�U7,�e՟lRtf|��\O+2j����w�H�m'�6	j���,���v�{(��9ˤ�>��2߅#��L��Z�\m�@67�hZ��:x~(
�"���u�D�FCaNC�cOU���!���-�.�5^�ޫQ�ه6�{+�����������85
	x��^���w6~��k�E
P�o}��޺ʮO�! �p��c��^�G���?m7=������E?��L�W�u������`�VphZv&����u=4n�k�.*�3o?�bu�W�Ifj�D�mQm�8���G�r,���m�bsq�]�}���) ��e�V�co5{��az����<"3�|�����I�h�u�r��MG�M���&���J����o��VY@B���Iij*_{��^���-�������u:x�L��zu '�H�[�Q��"�D�������@��l�>!W�3f����u���u���wF�����8��R�J�ψ��	�pɳa���Sڑ�4��ŢR�����P��N�隂�y�gG����t�*��e�T�j�֛_g��	ў!�Tq���J$<�K�d����!�H˩�b�8� /;�k<E"�^ck��xN���$�zF�ev���	�"Kk��ʏ�o;����O��{�W/q�����
X#b]
��&5lŅ��Txr1�V���'�1��y ��j8�w#劊eV��1l�>��K|1pw��+�e�1���4Y����V@���u�!��(U�nܶ܊��jgS۴mCULy��:�\��nql��{���0�$nd�|�aћ5�*�_�V�jE"��{�����+H�)@���$(\�9�e�m�/I���1T`�>������L7�9l�PE B|XF�Sc��K�w����~l����e� �(8�v(ɨz���O|�o^z��`t�}O?���C�K�x�4�������,�Gh�k�8�s�����i�Б��$���p*���l2��
�j�+o����S{ߵnqd��z�Iԓ]ج��ѡo���N��8*̛:.391�rZS����@�� ��N�`+����\.P�\Q���2IW�M�b�����H=��SE���cL�϶P��ܫ��f�~;�;��©�����Tm]�����!PR�~ۆ��$��O;���+��z���I�Y��0R�ދC:��-M�R���=�w�	����6bN����b��4��W���T��(��Z$
��1N;$Y׃�*�d����F�B��q�g ��[v�Y?�h?c���I�=�B%4�]���wG�����(��>K��h�N��'�^�a�.���x�8Z�))�n�>X��U�0�ާZfQv�'�1Q���q		�sÀ~P� P�S0/���v��4��C�&U</A�^���eh3n�S�6�X�'�IO���!U>���?<��/�����I|L-��}��L5x�$��M83>>+���������8� �� �����%r#��d%���/@Ծ�θ~mf��XwD
����Z�� ��O~��2KO�X5s�|(Fo�z��3��K���f/��$�����Ũ������E\~���h��P	rY�k���;	�i�#jI�1�Ш���C=wB"c
>�ϗ�:jwd%�#��r���Ygki�
J�!2��>��ɫ׈x��,(�T<�Z���8Sj�qӓ�7�=<�Ka<b7��G��lf�[V��4�e]�y��F?V�@�vv�PL1?xW�^H`�p|@,���e���"�o�e��b7����?9"��;�xm��/��8���kx��T�G}���ڂ�r�'
ajh{��b:���l<����5�r����{$,1#�������O���j�nU�a*���C�
�t	0�1��/����.� N����Q.o|������JR�bfa�]��¹|�'R9s���7���8�L������'3�a3ڄ���za/x��̵�aD��^< ���_IȖ7��Mu���~d/��'�����\�\��ʁz���E8_��FS��\�s�A�j·o٭U��I%�(��/4GB�\���:����yښǖ���2�08(�/��V�����Z�ۏ!^�Ea����%��q���1W�l�է�0T;��eS1���:IP ;������^<���EJs|Bw&bn����p�UO(j�!�ST��8�Kb�m��=�+���rR�:���2L�ӍJ_W��}e�4��͓�G�}°��?��*:�{f������7c�n���W>o�!�;`�Y0��� #�l�*(�ف@� �`�2}�!��q��9ؽR�o��?e���<���h��������$Wܭ.��H��̂�`�Cbj�\�����(s�IԿk~@f������[�j�^CA�:Б3���  m�HL�^y� Q�!�z��〃:)�>�)�C���Hhx/Eq��0%Ro���t-�khM�����;�@a�{r�s� �d�5�{�6@6ۜ*���L���\�1��7F�w�rs9�N%���.�#pC��`f�s�l�@��g`of�#�����\��n!�k�D�H5-��*W\��q�ɜ�(T���Q:�Oa��">���[4tO6�MϫIK&�F���*�yvӍ/D���F	�.�ǰ�M)a�  �:�ⷶ��& ���~��ZGͱ�"�V���T#�$�Q��NBf�A��y�o`�����kQ�j$�
l�?P.M�