XlxV64EB    8af6    1f50saf9����	������3頡z�Ro�x��,M0"h�ݝKYR��>�C�ǎ ��鞖�+�ы��h��(��M�a,ݣ���� Y �-8���/����pDs]>i�5�e�
{O3v�Y��]��7��x�Ql^5sx6�� $x��v2&s���Ob<Q�,��q<Bg�V�5����8�	~�S���w����h�L�":#ǫ5�z\~�?$44/�x+�`�����*e�͗d�J�(�L"#,8�:.6���oP��E6�Y��?��6VB!X��'�;ࡨ��و><��y	�4�����������͈�6�͋�M/�ٜI[*�u�id(y~�L}T�9�qMܶx�1��������H�f����$ ~?Ik��O+Xh�QU�X��ϡ� �#κ�H��jX;+�Zt	4� ���/�l��x���z�B�ќ�;��+9�2�9IB
���$,3�o��s{�'p}�[}Ӛ=�v�hJ0��6(Ɂ��u�F��A���\'Ʀ�`����L�sk��ֿ�l�ZF�O�H�X��xگ(�{��uF(� �~�XnY���WҴ�r�8;W�t3=��s����`��s�s0lR�k/-�8�	��h�H����YS�9W��:�'o���\��(�f��ve0b�d�c������ ���GV'2���� ������>���ͦC�����ƪ�n�c�����m�E�)��T���P!��"���˴�)�`RӞ��T���؄��B��M����O�h���:��!�zm��x��_�>�[
J-�l���d�v8?������u����b���@�B�g�~����?[r�@k"�uQIY�����1���*�5^����)��Ko��lOvfj�7�X���l �<OV�6⯇&Z�qH�Oe�;9�V5ј�t����Ȝw�2�,�p�݆F��_:��ӗ�����o*tM��H��`:� =�6�Ñen!�2/��>l�:�ƺs���}2F\����25s�^11�b���a&��4�x��q��G�q����>@Fs{OY>��Cj�����G��B-�Ƨ1�^!܂�n��3�x΋��O��,�1ZC��t&s'�n��:5�UƊ����9P�E)����a��K����r�n�d�d�~�9[�}ճ+i��j�c�� }�nW��������u�e��sg`4U"�?����܉ o��̀av!߯B�������+��v�BJ�V��u��B�o��j���p��(g������? �|Z�i/P�9���Z������y@�`ʛ�Z���sK�<��
�+X@&�~�$�l���� ��ˁ<�_�����m��В�sr������������[���&����{�=�/��d����$V?x�1��y�a������������hN+�'�P�Dԥ�A�p�ho�� �\F�f���K���ÕH�h�T(�ADx:��C��`̫A�X"e�;'FC�}��u�u=��WU�w���^Q���hB�ɍ�ƅnK@R6���|8RBi�������Ȅ�eO�������ʔR�R4ھH�X�KZ�6d����)�
�_���m�ZF����j��U�p����7��9�YԲ$_����3$}���3���q-�:�Ye�g/�.KRr׫'@��� ������[C����G9��mV�ܫ��P鐫��Ԁ>b��˵�.���7��v�vrh@14�a���F�l��UR6-<���/��_Z�2���E�H�C_�K�_4Pvg^ڶ5Dp1�q_oج7)hV�hM��@\����?�w����P�C�T�w�J���w�J9��$�x�<o�)�n�{U]�Q�[W~Q�̨��]��i�����@��'��Ϩ�9:~�/#�/?��!��.���j� �}�L��t���
�u��)&�A
���ڕ�,�1��?̰AZ�j"�N�f|5`�JEV�|�Q��z7�8����6��q�V�e��Ia�N�qr���<�}�<��Wf ل4��p����OC���{6�e M�e�tV���E�z41<�RN�����q�%nӴ��H@Lg�4��o��تT#+�|ρM��;�׎�$<}�<�%O���*(�;{7Q?��n �?"�hie�R���� =+�ku.68�@U����&O�ݕK不�1���e��Ձ��G͡�ȥ:\�ciw���<lD��C?�d�����c�������{M�b֧��,,`Ϟ�%ͤ�:��+��)�e��`ԧ˴�b�ؼ^7aե\������
Ě�F/n嵕md{�X�f�V�	���l�+;�M+��l�����/ۦ[0��Ds��	����<���(o�ӓfd��㸖Q�#�[�H2��I��KR�P����e��(E��)6����Ы��y��Ã��*��˄��_����� �N�"[���� ��l��`9lM����3�@����EbA�*Ml���q!>�#�"p>l�fM�]`�$˄��3�[S�*��$i�1����~�+�<��c���=��ّ��V�u\6����L:M����`j��c "�Q�%�	�l���I�n�N�kM�`e(��k]x�	=&"�=�����`߂�GF�l����B�囧�қ��X�sI=�� ����Ă(i�''�S����`zX�zĹ`9ä�ᑆ�{C_�W���;��������f��PP�3��e!���� � \�����s��L��JcȀQJ��x��A� �}��v��anly2�*�� �x�3�-�9��)Vy�J��Z��d/���V�H�����J�ݻ�J�,a%�]&�2*���3q�sL�Ĵ;S������&q��+��8�`�D�w�(q1��I�|C03��[՞�5D�D����x61�Eb�m���x���<dNE#E�:A��®��ɍ헾̛3)�o����2�*�cUhs��]�oNir�%���M:<��>:t�:��Jk�I�@t�����8?zc��,�X�G���n=Qƿ���hu	�=VFtG��G1F�Φ@�S�N,�J�N���"u2ņ�L��z��&Q��S�{|,Mc�4����`=���}'S�G�����3]�:�I���87�禭�B��	H�T���Rm�Q���6�m�s,z]�#�1�$�;�yF���;ի�{��ԓW$i�}n^D�6L��U��1i�������--L">�#<���a��ȁ>����<�������cz}Q��&P�����o���1�T|��NU����,X-{��JA��p �&�E�13�L���q�rzR�I�w����T8�ō�8D@8�r�>l�X����� �e���0Fz؄I�Є� K^[�8 �
�&Sf������.��>�7J U�;XҺT�� /�]L���p��C}\�u�fA~1����Ϡ����>+p>�I8��B�r��W��N�@9��i���l����>b�t�������N�rNM�ՠm��j*f�fX�'QpF|X�`P,�bg �ԫo�% ���/���3�V^�3"Z��D䎂�*O��D��"=3ҶBR!|?��k��e�F���IBء5���Qc�3�*/��v6 ��V,TP���&��݃%�u#?0(_a�kG5뎸�Ѱ�A(��=Wį���H�������Jy�Kc ��ް@V��������)Jҋ@���_}:3�����>�znF�5���D��}�Æ����>��4�t���d�`�ǥE���6��^D|}/yM׫^�S�[������������b�j�ҷ���0I,�f׈�`v+��͕zM���TI=G��-�����|�n�K��,t3��=�m����i�mĚ��W�� $4-*p�{%�����oh4�򊂑�)��q�=7ٳi7�I4�H�?q��A��3Ȼ��|}��P���h��2�=VUw��4��~��'a�їE�-��L��]
�4��f���!:��g�i�Yr�$A��?�QG�*Q%fş�Xs4�e.deN���]�`p��0O<��G�{3w�����7��s�n��������~��[S�c�r%'?�S'���הc���cd�t���t��f�3q���2�a�� Za�yw艥�X�6�7uFH�Y�3*�Ҽx�AG*���}d�h7w(�y�}-��i{�R�"�y�:����N��K�{[E"��@����2�z3*x�,fru�14��?X,b����$�(��`u�;RtC���$��G�2D��k���}r��xxtJ����q{��������(�vXv�6����K$�;\B>މK�%
��e]�c�)����V��2t!²/��-be�V9��-oV��u��a���W�0�/��Q�Lg*��<�����ܒg6V����MA�|O�.R�#M�JN8y�7y^���5�ז�xu�c7P��=�� c����%�K�z�ʣ@�s �6J͊`���a�B�����?�T��N��jý��p�m���q��$vP��꧜/�d���hk�?o?��z���*s�l,a�&��|�t[S����w�]0\r��H�������dnBA�I�oX�#�#��g�;�?���M1�2��_�F��.��9Pc1����{���^^�XL�h���gO��1��9������7��vd�/�h\ށ�n�H�xY\���ѝM�-��<Z�C�i9����V��N̺�t�],;'P�w����*G����E�k�1O�\E��C�ct�@�.�XO�k/k��j-\u����:zpa��fxm�E:x񙴍��|���C˖��H�:�I��MA�d#:/��{�f�+�ޕ?�?�q�H�I����Sɂ"u�J���SyP��nN#�~�_-��oē���𱚆�����>u����N&�2^��j"�ӻ6�3������M]1C@�rM��]��,w�3�(  ��o,!P=Y]��(i��X1/k��h�f}�[���D�U�sn��
KC|x�f����cEۙH�\u]~��$�ڿ��ݞe'�n_E�73��R?��1J�=)c�4 b9�JQ+lS� G]�.�����c^:K��;��M��]O��Fb��,�;������'��#Xx�)w>��-���{��̔����K��tƦ�9s�^Df1WqG�UE�֨�^��GetD*B�5o�ޒ���qtǱ�ao�+0��i�R6@�� ?h�l"#�h����D,��+�52�?r��L���P��0&�o0yv��Q���t�nY�G������<W�b2��"���-�=(x� =�K������/̝�0�gt������m�&�<�.�	+yE�U��؝�!��՝g^y�3�+��d(W�pW�ٮo.|C� �aD�ӄH�� �'�{�}�&U>q.-�_�K�� d���>��9��Nt&��Z#w��T��i�u���ld���Q /ȮE9��ӽj��h�L<M��OS1�a�+�E���/n�L��%
�t���;�D�ɽ�������\
5ӓ��b�{2�L�F6�d���Hb��Qm�؛}o�xp�!\G��ӣ$�X,,k�.+l	+�Ҋ�AK�8V٢�	7ΓZ�{=�9�c�Jw�
��~��D0�o��A�<M0�z Bs(4�P�5�R�L�D8��\3��Vš�I5����z�d�O��V�!��a�~�O� (�@f3\�!��)��g�RJ�������r�[S��R\�9>*,����F���u�&0������ ��E��,lE� ���[Rp�r!��׍U�Б�灙>Y�%+��#Wk1��O-1
���Ԑs|²�=�qܨ)�I8�Hݯ��&M5U��������j��\����U�9��k���v`��~kY����&?��a,Zo�ߌ�?Fq_3I��LVS�na����6;��ɖ�<�)=~!���t5���l�+��,,�{����X\[��y��Y��0G�~�Gd,��z��6�io����5ؗk𗒶9��>i����9���$-� B���$Cfa��ǟ�>�+`A]�*t��_�}{��Ă����(U�#�u�?I��D}9��Y�7+K1P�MZ� '<�S����n@�$�μF�������}�������3��Lמe�E��a��['Z�:�Wu �R���@G���䩡x��>�q�)�1櫳��I*Y2��P�ߥ���Gp�c�Ķ,�UR6!��a�=�G=�פ\���يF���|q�Jd�3�����6��N�A�Sq���]7�q܉�����@ێ�.q��ӉQ���);��4f�X�q����D8h�r="<i�Ea���}�5i�hxVH!v���8��Ȝ4t�7HĶ/:A�]$�L����7fp��C��%�fs*'�^�|�p9�ϩ��谘���+箂�+��V�9�W3��N�k���x/c��^<�a4w��������+՝�k��Y�vm!�y�r�Fɚ�����>��].����Wj�y�N$lIM�@0B�5+u���Ʋ^byO*��+>�����xS8�mͰc��q,�i!:{�ƒ�n� 7������b�g�c`�O;]�e�hLa]����BgK�^�6-r��lН&�v�K��R���)"��%��a�y1������%;�+�
v ��L�����y_c�i�=n����v�8,y��Po�Z��,�'j�Y(o�����Wd!���]0�o�=+��gq��՟���J*�a�+�j�����9��l�^�9��ٖ(诉C�:���h���![�I%݅"�qj�
��¿��k;�Uk����f�8,�戼�-�W�=�w���+u9U4�Z����.��jzR�0 ��bQ����Yt�wZ�/P���쪦8�G7,����\�}���1���'c�U��NC%�J5��/�����q2c'ܸZ��v>�wE ������Jw��7�lF#��w������r0�4�%���4�k{�ܽk^W!�T��[ډ8�1��b���D�m�yX�狐z
���✤������Kydh���C��8I��P�2��B �T����Xes��BKm����u�/�a�ֆL`�*-H��G�c	�f,@�5����W�����j)fla%�qE�K5^`n��)uo�#��$��چ~��c8?q��"��P��i�:Q4 �	.hu~$�����cz��)!��Ч-�A�8��5/]�~�x?��UzwR�����H�y��:��|֭�&��^KOUU�Lp^�n�����ʄ%+
l�ѣ=|q��A�I�� 0twx����Ơ�R+]��]�yLfytk�,���l�A��z�6P�r���4���Ȩ��\�y�8H�����y��n�5�����$-�gU��e*٪�p���t�t�?+R��^i@e�_�/�HN7U b�t��N�c�U���X)|�N;�Z"�V��7+�/8��w c��h��:u�0{��S�~���c@:F�S.�ت�琯�k�rt��=�T|[��5D������d�Uu`"U�dL��VKV�I���BE6 ����`S~.�l���_�B1p�[��l�B=��)�ix7i-����BTݺ�:��������a�
�s �x�xg�s%;��Am�UW��0��a^���E��[��F
\��мV����F�O��w?��T�i|Y�%!-U�Y7I�sU��x��`}pD���hՃ��[�N��lK�&��9*-`��1z�6�o^��f�̢2�=��m�F:���M����i�d���&�/�O ���e����D��"t�K�lLӈ"V�C��g�i���J���.Eyٝ��O˧��XyX�pgbl��P��N9