XlxV64EB    1dfe     9f0��P�C'��b[��}��r�Ԝ���|6vH��"R�1��o��T����agUIy[�)d;�}%g�x�t�x�bhh�gj`�Q��Zy<�?_IIcm��<��(����?Qɻ��-�󋮀��sU�R@B�N�
IZ|5��0D�:X���_�.rd��@�T�&�������ͬ +C���u�KR.��%�~p�R��&ēpѧ|m�â#P����=0{�P+��O�������f��^PJ�MV�x�����V�ƞ�3b��J���@Nh4Bak��E`��JSu�@�C �8d�E�p{V&�]�i@��9�h� �P`��xB�q��O|��j����d���CsCהi�ث��n2�T�!�iX�c��
O�Ѧ��(���1�k� �R�lb��8�g��L�3%8�f]tW�~��ۢ�}E9bk�����z�sMh
M���f)�*q��
|z��Q2��&3�HS��W�vP��Bf8Oc�a[�G�Y��=�b6D6D���Ⱦ���:Hzq��ˡl�(S�7������� �<�|���I4H[�� J�e@g�&���@-�-��a��T��|������d���x�8����І�1%}D��t3�c)��p:���;�:���y�����!�'���J��\��s�i��LCnj���JKA)��$�����:,ԹSt][��)ĺJ�$��o�����c.�-Gf_T���e���N%	�֚�(�*�F�1Yl=fT 撃W ���IW���F��R�a��B5Tf��z)�@W,P�Œ|�e�m]!pT����y[XF���q1м�gG���)�}���,(_�x84� �H	�O�^uW�m}�9)w��̬�S��S�,���Q�8�x���g5��(TK�
�!���|�U���e�λO�@؆����_���h�J+D�.7x�]N9\��B)��Å:I�b�ѝ��h�Y���WO3��1�پ匔t��<�n�ݾ��kg,~�y/�W�-�D��=��ŧ�1�3�Y��	�]�g�tή����@y#n�?[׷+̈́�x����HWQ��e
4�d�tے������ޘ��)fLb�)��w#4w��0Ŵn<$f���E�v;�Q5���ԜK׃��?0���gU�*�X��@���~""s�����2H��am���>8�%�u�,Q�vze�?�������Pn���<j������@�!�e�8E�c^�4��f���f;����$ﯲ�Z�������]݆���sO�p4l-��>�
O��z�4�+�pp���D;��{��zZ�8?Šp)m	L�=u�)^�W��v����ڍ�؝����]�S�Gy&٤1���fM�9���=*�Zr�	R�QI����AAq�4N-fXe���Q5�5�(���h�^�>�(�C^S�o~���C[�d3�3H����2�����L�	�{�;��kA�Tv(`����a��㟾)�H�c��as\V��T$�X�2��X;|�iS�3�:Vi��z�Z���N�ֻ������Bp�M����P�z<�NT3�
��-,U��>	��Ŵ�C��߶�-�#�JO+�dF�/`�X���Ou#�]`��r��Z�VO����sf��k�X��)F<��7�0�!^���"/9���~�,����~�:��<�13�Z�!��Ad �	��G7i9�r��A���<�%�� ��&1-]���>?I�k+�Qt����t;Q9�P�[�5��B����Sފ������7�K�R�sR��/��n1�Uh�@s�tY4s��=��؂��x��j��D����Ѷۉtc��^�&&��VJ\qX/���1YA���d*!7�țO�<9y4���smN���ܵ�#�4~}}y��!��2?d��>�U�ך3�j�P����ӧ༠�ר�bk�Y�/�(�T�ݣ_�`ϕ�n[�0�i������^���S��K�ӊ�W ,�#\�W;3���w�	��Iȫi�v������eo5KlU����`�9�/
�B��{`~��X��w&5�L�E��o4!8��bv
5���$7�U�q�ɝPp8<�� ǚ�:��GŹ8���D���L�*���z`U^9l��UvAlK�!���B@> ��5�:%Ş��K�	�tD��|_�2�{��{o7kU��{�r���Ĉ�;��E���J�$ϛ�%(���ئ��=�Y�[( j���g\s��f"�zޅ�(A�JP���"O'�н�m���������Us��OZ�#c�+"�y�n:� ��>����6նCS�"��ŋ�̻TO���`"]mǭ�Е���$0Z�BL?��kSIX�B";���x��Z'�"-��v��.��#�8"&�� �
��X�\Un��\�?kr�q��TX�⥿�WN�-��Bs��[�>����ˤt+���?_���p��Y84Y�|197aƢ�GQ�U!6��(�7�5^�����fD�@�+�u<_�`^H8