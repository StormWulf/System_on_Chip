XlxV64EB    237d     bc0�����jg��[џG=3˂���J����0���"���6/��Oc��	��������f���Gn5�WnF4��ss q�)=8jTvN8%��%AXlЙHz�M���22%q�<n4��Z0� �(:��OWV����Z�(A,<)�P�UQN���cL�ʫc5�R��&���;(�!$�D�`�=]�_����A*�x@��዁�����<8 $u��s���O�j�>�A�#��]�dC\�3��$n�T4b,>2�k2(цu��4~�D�G�}Cm���Ѷ_����t_b�I�f1�L���𦼔d�=~#����ʷ�Ζ"�}j��IL����& �����FA2�T� $4׎�i,M��8����RS�_i�/=	�שq���Sg3u8|�7��WmG�=F�@��<�oy��,�oP��f��7�\9��
�UL8�-�1:K��I��S��(#/XkW@.8)`W�/���>�dǱ�0��Ƞ�mO�0��~?�QX�ߧ(ݎ��o�Ԝ>F^�>�8Za����m�3��L' WQM�'"F��������Y��Y��������p&-��xu����l �;����5�����MY�3Ya<!�����U���޻���S8�"��2�J�[�Ş�7�nr <����cG����6�ɗS�Ç�]��.��b�YmE��E�E�1�}�Fg#�S~�}�Vm�������"|�!��&-��G#��[�vo ���'Xp+�ݒ��WL�B�����2�@�t�@a�d.�&��s0�Q�xC?�r٫�A���ie���)4dM�_-T�s��|�C���Z"�)Y6�GK+��z��=���'q���^8�d6f�&��������pr�l�rθq¸��7�.��Q��p�����q=�#��T�w@g_���� J����Ċ��{PU�R����.�%u�Z��Qg �<�����>�����O�dQ�tlᬨ�*Z,gC�i�OKE���$�q07��-�Y����([�k�0k��[3�폍��Z��U��SUC[�{Y�s�b\�а��������U��ά��U,'�	�8�6���F����c�|�-U!�1�W��j�T&�:�|�}�j�<fa��Ĵ����H#>�9���s47�A�a`�a�>?�x�,;2��yc��U^%���8�.�RAªx<ni��ˉ�P[��T�\������V˝�O$��&�,�_�%�c�Z�8�ʞa����g���n�[c�8�3�2��8�Bl�j#��� �[*�zB\T����^�B(y}�jc��$;���
�A��tԳ�	e���|i�F��6���Zj^`�텑|g���탑���:_���`I�G��~ƺSn�a�X��ȳ�z�X�Zݴ���_��0IW/�u��.Z�.k�Uzcq�P,��)�$�@�$h5�lG���oR��%7.{�F�z���=&ym�B'�)Z�Qa�J��_o�q�,$��fFQ8��vt�x�B�=�,��-W?�?� �V|��w��vie�-���9tx<��YO��EՐ1骰����Wt:��0��-��Twj�	^d��d�!���9ѧ�	רw�0ג`g�Y�V5N�J�2�J�D�\w�@��0�Ԗ��R�0]/j��Տ�8�7�r�v�m�t,pv5ߛ�d民���r�M5}�I��-�eKG=��b��Gb�4 QR��rV�ki��x���}�v�G��|��/u4�U#!���/$��q/�u��Gv�3 ��3_(}�o�4��n�]*�C�m���]FU��q�%�or�>����Rm�7����(��:*9���@�n��*o�U�	�rH`��â��͛��<U��B���cy�Ԕ�LE����gPA���	�yT�=�V�ҀI�cfe�w@k,+�h}VJp��\{\4{_�����g�*�dic��S��/ӘRߒ�}W�:w+Ǧ߼�#.�;����2�DSս�)�KN/�d*|pc�ydk1����H��@�L��k��-�$��Լp�ci����IͲoo��g�)&�0�
R��g׷�l<��@�����D��䦎G���Y���YN�-�t i�"J[�K���k���"��s2�����`܈I4\������c?��
?\|3wq��!7=Bj�jOv�����0�|��jb�j���Cv����ۯD��Sg�����`�R!$��}��|��DZ����?�1]�$X���(h�N���gq��nP��)�=XAm���Eظw�Ҫ^��:��d��AI�]���kT{�m�u�<>�n�:?2w�s�h����c�#_]>c@�1�p��R �5;9�ĸ�R���� � V��=r��e�����]=A�����i΍Rl+n��'�4sR_p_�1�#��vֽ
>��Wb���>Y�G� ���w,�sԱ�2��a@!@$C��o�}���˖8�\�ƍL{}���3i�)�|n˃A��`�S�T����6=9��m\O{���1k��6t��a�����NQB;P��P�'�x�	�O�'qpE��x5��M��
u�%��.����ZUm2s����)H���v>g�����g�m�BD����]qI�YÕ;���u�[I��A�λ�?��
6pI�����@�bfe�r��p�����a	��a�R���=kL8���M�ˆ���ޛ�O������\G"Ҝ�P�)ZvqH҆�7�=����dƂ��8$���v"˖%	z�0
�.�Ŋ�Z��(�[C}Sd;N�V�F�$)�#b��kv�aHV���ha�0

ͻ�#E~�� �tz�a��+%/�%��g�r�S8��o�p���rѩ!<�*,b�-��Y��_�c�wP"�EU�<�{P�r]3I��~�5����+M�y����g�Y��mU>��u����E������ۮ7@˖Jt�Ü/,�o^Rb��g�BW��{R3{���� `�"���