XlxV64EB    26e4     ba0$�ʖ���Z����>���#�Ʊ��D�2ւ�-�����.I9�� ��*�R���M��sZ �ͷ�7�2¸i���}���܆=_�:;U����S?v!5���w͋��4kQ8�S�h�ns�Ϸ���d	�����"�e
hC�7�*�cpEh���I��^�ʮ��:�-�� o[���>	n��]��,r��e�|DB0ꑙX�t=�S����XT�v}�po�^inK�0;=_��3�C�۔�}?`��Vp��9U&O���R�e���9���������������Q�~Uk:Nr���)� ׈mIU�q(3�?�����uv��;u�`�jJ<<pQ�,�;@��y}�3��3�G;�X�Ao&�W�|!�	8��^���� #gh��}ֱe~�s��hm�wU�T_� &����7��! &.��	�i�<���	���~��/����Bw����`E�%�Y����Nk��yU)�d_N;������}����y�#v�ğ�y��G���fcAwk-����B'�w>�/��KG�Y<}�aم	�a	2Յ��gΧ�K��-+�\�߷ҚW��3�}Y��m��J��Nf�����iR���\M�Ϋ�Et4��	�$���00�SYV��@ϵ.w{-��u��h�Z�Q�.�k��	��d;b��Ā�9M��.2�ܺ����t��cY���G�3O�_W�-�&���['ܾ�D�k��lVEƁ��pO����k�:�٭�������v�
���՜�'j����*I�C�|��w���'�J;�8�w�ɎѲ���:��_
��:�6��?�R�Q��F% _�32����K��,D}�v�P�.�+p~�(����׫B�8��`�L��t8�3��<��Q_l��.	����k���|�2�@���k���ʤ��o �����@J7TӦ)s�QT]�֥nz���|s����@�R綃�
��i�͕�24�!���Tۆ��`
��\N��s-�ţ�c��$;�<���d^�t$��r=���T �Q��6j���I�����z5�_R%���pu�s��<��!��x��݊%&�i��(����{E�S�߱u�=L����Ğ�&�����.�s�5A]̚&��L�0������_F��2:��W��p�/ �pd�y|��ڢ��VF�HX�e	z�D��Px�bɫz\���|&��ȣ����|3>X�~��L���d9Q}�B�-%��sԻ��fYi �O���~�:�$x���p@�����*8��B$'����U�@-�(W�20��n���|�L\�P�gL��W�iGT�\��DO>)��D�_:S�ni�~]�k��(�>�vA��o�O���7��PNr�Z;m�ʋ����	�Ɇ��d�g���^B���� ����rO��I���d{�29�"���I矾p�_yEdSޢ�~v�T��-���6[�Y�� �Z��D�K�$�"����k�����X7�����Ȋ:�p��RsM�3�O��a�SO3��l;ϼ&E�,�DA�c����iYb-"��Xi�>8��7�Q\��y�,�Z�ޟHڪ�U�	j�]�z(�zd��ّJ$��7y���ns���D�+�����w�k��er��72��� &tci-�\|˅\ұ֪@�'��5:�A R��p���&{y�|���ҁG%�R�%�FJ4��G�J;�ы���<R����&�oX�ڏ$�9�T�꒏��t��+֌z IW�ȡ	�g	h��Jq�fTUC�:�'�K��b$��c���G(�?�S���	��`G{�C��
�nyx�r(R���,q���K���}$�e��[k�]0�bI�g��g4���	�:�6�������R��8���MCܶ�q=`�b1���:�'�T_��qP�ߟ���ć�ɵ�Ջ:��5�Ԥ{�Wn�W&H��1�u���`�X�d�^�"g4>��ki��R$���RU�5?��є�s���'����/ڏ��*�|O���	�q�&�A�W�������`�����)��Y��^��R�[m��A�'by ����,�x�urD��<Jk-u�"�V*x�C�F�(p���w���a�ѵ��G�^R;{�<ttn��" dƟ�'�^�M�
�4��7��g�3ٺ�HB�0�tӿ�>%6���&��9m���������A��P�^'�����O�U.-�����[��̅8��h�g6|��[]4"g��`�U�f�S�Qe�5,A1J�����*-^�{�{ʢ��*�w,�}s˂JA��p�B�v�d���b�,���g�Ź�����%�3@#����1UcZ�ٓ��0��-Qf��	�S.��8,l�"�+����0��m�����<������=��bb������O�~,e�3��g����+�s�_��d�K��S�9]�s�a���!���]Q�"�a���G�ԡ!�B�@qt����G��B�hCף}��Q�z�i�j��%{ _��В���*��a-��v�"�vQXE91�[�}�]@n�_?�ݵ�]v�б؛�)覅6���ߊ�������5zn��f{B�{��i@l��/����ꩍ	�"��R��[�����*�#�麞�=>k��[�k;�C�c�.�E�����jG�_��.��J���7Q�i��<�f���^*�M���u0j)ȳq��$D[zĳ���D�,ޗ[,�f9�qO�1��X�Ee�3|(�^#�iu���*�Mb�����+?�������[����EUD�h��#UV^�~��H�᭔!|̾�?�<� �:�5�A�����A�I��N��H��� �ԣ�_q�����Fwó7G�W;z��'5��i�����#�>e6B²����E{��$�s��ڔBZ�=B"�>�������TU��B�䛌�z�T