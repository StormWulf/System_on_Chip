XlxV64EB    5cba    1430%����g?���
����?��l��D�����)_\�y�}��{xv���Ss�#��?�ى���f b撄�T���N�Jv׍��m��S�6Z�"���Ie\:�s�ý�hj8�K��F)C�7�pE��\��o������T�&�ԣ"}I��y�6+�����4�d=@(�dCC���I������[�`]4e2��Ai���hh���b�%�iئ`ݮp��������=��|�rVL�jP��<nA�{�=̨��oh�e��"��
��b�����T�����h'�Wn^�㳸_"*aP�"8�T���_Xg��JP^�b����)�`Nޖ���U�^W�^AyJƳ�l�|�cA3L�Rc)����f�b`ܶb��=�< T" =����~wtL�`$I�&��}2eLf
.��_ƧՉjj�U�ǲt���(2���J�wVٝ�cG��8w"�\Yn�r]�8x��FBꥁ�"�;h�-K��s�����Ֆ���$Q0-����'ӧX��f�@z�]0�אQ� �{�Yg����J�&���z�b\K2c�<�*�;������DδN�ޓv�x��n6�<�"~~jy��2�e����<I��sh��+-�0�ʵA��
��E�.��\'��8F��+���7��
[�s�~�$z-�/����+,������6h\����?�q}p�Zv��{��5���y���d�v���������!�sII?��b��Sh�x�~hտ�џ� ����� �
&�pZ�t�W���?����mw�c�'�Cf_�r=��#%���q�瘠h,ɪ��Ť�� �a��~��IIW�Va�\3�\��Tw��"ښЁ0�q��K��
;Dn"̀�}Cu!����jx�K��N����4�*q����9�Td4�}؊e���hZ,/�|Sog"���ď ǆ2�1�6�=!�5��d��#a%��gmO
Ղ�U[;�iԾ4{!��T��?si�D�t�/%�i��[�XW\���ds=�H�*�x��H�,Xf,9�i�"|��==ǥ>W+˪��_ ��U9�å �Bʤ;�l��a�����Lc�9W�};Z��7��^�V��9�톟��]�o�2J ��8�B1+�iQǉ�5~B�5=�.W����v$�"�Y+���tA���j�y�p������p�/䧬{c�}���%��X{��e�tD�DFr�f��F�(���BGtꯕ��š�T�r_v-{%l�Ve����!r��1v��W��q�1���j5>J�e�U$�2~�����E^j}v��a�v�*�kA�R(�g�^V�q��\4"�T�><����J+	k�Ɨ��n���n@���M��I��a��F��GlN��-���	�QL�o�C@؄�n2�%�U�1�_.��ڥLyx�R�wGԏ��v��-��qe9����64��ף�+�^�O������74�������%�ק�݀đ��m�A�p�6[-C�N��E�E`(�+�'1��08g���[�Ұn���rG(X%�Ӗ7(ߵ��9U�����e�l�ϻ�tv����"��q�����:ř�/���z��)���I~9�.��]��!H����
\���ti m��l���I��z+g����Y(=��=�ƅV`@.�5N#�Jyk�h�}���W��:�:�������> �U�@EZ��#/:!��~F/L��c���d&�w��
��r�C�pNW�������Z�H��U7Q�A���������ၽ?�5�H~��� 0�k8f�[���0�xu����۶����g�>Vߖx��y��D�d����m[�Gu�V����j0v�����|OF�o����Vmd�3�WM(ղ-ro�����?j׷�/��qo�H�G�ޚ���˼�7�A7����K�T!FJ��*`�1�P�`p��B)���Cw5���	��dLÆ��ݗ�4���Y��H�T�A�"4���|nUZ�
���71]
[3�b�b��qd<�&ܠ�t�d���f���D���y?f?�=-ўh�	
�/rh��bm��Z�����zp�"mׄ��ߝ����g���������t���O9��7�d�U��(	�>�m�S��Z�������vw�TT'M4����M`yȈ0�p��T��u(�Ә�g��ژ+m�
�Y89�梵K}Y��QP��X���1S ���3Xb?�D\�X`�e��&����͜����+�������%g��h��%��B�C�z�@��+�x��^�5�5�A��SP3K##+{�c�-$?!�ܯU&-l��VrD�̋�**oo�K�A-�� ��>Zqȕ�t�i)έ_]�ݬ�>�P�J����]�s%:�����K�&F���tq6a�U#�xl�a�U�ǃ��ʊ�Y��m���}M�������F[A ����*��N�MR��)���_���Y�	���؞=Y�韟����c���>6,�$�@naZ�#�WA$�=���n�E�����-���R��(���J�%C� ��,���v��Z��T$ߵ�̴(���?�}g4WU:?g�,k��W�{/z��뿦X����=K�тd�Z��Q��W����k|��Ҋ����/Y��� ����aҾ��ػ��?M��BXA΄� ��=}�K݃���S2��lu�]���<{��'#����9��ҁ_=Ny)e�M�@[JS~��<��
�lX�;5�"���G28*�� s���b������j��[ڴ*?� hC�/m��j~ 
As<T�����"��X&��WL�у6U����7Z�P��U�S�x*�|:�Ė8Fxq�)�7�H�ٚ������c��^q0ەl�M�E���^#��N�X��p,�O�{��N8`BQCwbo+I�&��kC�W��u��ˠ�~��&ײ/�6لҞ�C�]�2=�"]��t��?z�+��C�IkC#����b��[M��T�q@㾖�>a� !��ubU6�G�Ӻ�땼�7����@Sh,����G��#�ۥC�W�-�ݫ��y7V�-�2�.R�a�(�RF�[�s3n�H��NaE��0�AkK�uu�H����i �.V|%�d��Ӎ%��h(��Bg���Swg,�3��79#��]�[��t�Rn�uyo�$�"�~z�������nbu�C�p�i�,��tS1:> j=��R�T�����8^��g���^Q:�AV5�����%��
8Q�..�<�dJ�NW�no+q6���O�K���.��Q�k�ʖ���jI��U��<��r�J��x�\�?�����̻� s4z߫�d��37f`��3P�ӵR%�r��-t��2���:萛��2�h#�`���׷(�p'߯86 �]�OV��\t�	t��"�b�2��6Vx���R]4o�Qg]�ȏ�̾r��z�pE�&��~��r0?�Hy>�$�$Ĝَ���e{ٻ�Te��H��H2.��p�d<�ҼW������=���q���Xu�{0�ƻD��N3k���J�2x���-�:�����W�ơ�bUӯKw�-ī�$x�6��E�E�� ��Am��3۹���T����NL`���{���dĻEP��J֩��J��5$�Ƅ*8��q �!?8~DpC���2>��M��&��nR���s�N<c�]/���뒉��a�{� ����E�"�7�Lբ�� ���^����"�+�H����̅�N��q&}��_bQ_X ����[��P���^&Q�T�$1-���;Zre���X��+��EC��RQ��;� �dsB��7�^�Y6QŢUB`W��&�W�]b~�F��Pv��$�*����ϲ#���5u�!���Z���q�z$x�c� @���"��	C촒$���%1���X(G������[1�+�>���D���f�}7D_9��eFˈݳ��Vu�*'���
�z�["�Ѝ�4Q;]��S. �4;8�����`^XF	,A-<RR������N���{>?�\��w��?������צ)�)���؈��"�;����/�\t*�\�d3�[��{;$���i��o��´Y&QHU��;{���	�EJ Hn�O���K��P��q/9�\A��Ⱦ�k��S��~�?9Ht�ABW`�)�>�o�W=�D��=3�F���j�u(���Z�'0Q�ܻ�kj����Y�ߚ�`z��LeA����ў�Z9���~��*4��j�d�2�aI��Z,kn3m&2����]_K�,ͨDI����n��iC
���8-�a��thFk��
%�i������:"�@���H J������+��9�h5��-��ǥ��n\
7?���4U���`�x��F<�êfVQHY�ō���+��{@�b"�"�4�7S%'�:�
�.x
Ơ̤�v�	� ��Pޡ�6�׬Um��k���C����A�VP�|OA	�T|+!S�q�w���D�H�1{qz�u�����tyەI�m�)���b��v@t1�I2]�N`<��R!���,�nl��M�*Nh;/�+�c|��:޶�V����߈ǻ
ҏKy�A~�6���fj�L<�G��cW<P]yw|��|ds�`:�����Sn���iz��QW�מ1�u�0����uy��-T���a�����	D�s8A,>O�Զfd�/@'ԸM3��қz˹1�~��P�Ϳ+��]C�OZ��j$兟C�I�����b|u�ʏm �#��'��@�9�,)��|����#�u���釋9�/�+nG��Wp���5���.6;��4��y��O2Vӻ~�N4܇�vM�� m/�94�3r�yy�(�e�"��u3R�����OaP��w�� XF�R�/�pЩ~�^��M	v�������xL `������kn_�����k�z�mnZ9L��7�hk�` |U|1�E���H
[L�m���x��!ě���j��,v�P���P�\Ř6H�Is���4��u��]�m繚���N8\5_�z���$�1E�����(:��_M@Xp�N�=�>���N�L?