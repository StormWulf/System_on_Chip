XlxV64EB    3eee     eb0q@��)��&L�9���yL�H���@�W0k���HN�zoa��@?tg�Ri} ����%gm��U�T-U޲�^�1-�#"�%yҙ���i�Ih�G�Zs3ߚ�H��4�s�,J���W \��u_�&�0�f�j��Ew�T'�_��Y�j\�e`�抨\w\?�tT�}���%&fut����5f�&���[���������X��e$H�E��ǖ�Z���P�l1�Y���H7��o�rD@���2����s���w�{a�T����ڭ��Ɉ�y��6E&L 9w ��A�fL㋠�������ʆ��m5���W�BL��X�\
�:\��,��T�x�����|ͤʜB�+x�Q����VE����<�W��,��'��Nk���;�<O+LS�C��	*�}��<�no�Rc��jF{�,�f�'SGg�Ty5�/��m�C&{#O�\7���q��'��*�^n����i�z�t�/���8�D�SK�s!����f2
sWGˇ
m���(����_
?qk��
n޿%���=�Ѡ!��s�T�d�L'D��z���O?�#p���R'��3t�S�Za	r�`_l�mۍ(az-ȶ�ߠ�}pr}yfdה�m���{��E���Q����˂�>��;���Q���\������8&�g�i�՟	?Ճd��'�kpj3��?\D��ћ���I뀍�������;��u�[�]���oc(�.#�s�+��Y[���-�Q@(Mz
dF�����$+��˘���)-O&����M&ѩl��t	]�X���Iq�4���mI�1p��030u�N p<�F�:~��-��v��N�B�I~I�%�����x��5Μ'f6Mu2���e6�����L����՞N�>������:�9�*=��[0��8��cYs����,ތ��������g����@�e�0�WMl�2"j��C$l�2��^���3��Yň���Q�0�x�t97�]�O��\�<	��9�@A��9�Ȁ��
�X�m�L��g6�3'n���iܯe�o�R�z$o�;�����0DU�e���>����^X_�^K��\��o�8�rm����Ҳ}7�-S}@��]2������gTDϣ�~QP���,{8�pFRQ��T����d(�ʶ��"���B�QWS����w$�� d�	�ʆ���u����U�A����b��,�o����p@y�F���^"��F^�P���?�<�4#S���f
`j�T��%A����2o�����[��<�nª��t�诂�U�z��2��pv\��e #������h����Q��ȥ}�y��VN���aN��
��]Z�V@3࡭8���n��ܱ7�����������d��D��.,�n�P_��Ӭ
�;1hos���$�;�Tg��j� ޛ����\�΅�S��P:�Q���_������(���#�G�ˣ�S��,��#��\1ǝ��ydS�:�v�D��h1;��*sm����?�X?9���n�x?��`��P��e\�1�ǌ�a����*O�O�(�������s荆@��>�|`a�#"D�CO$o8�2A�5�d|���W��o�-+�x7p�O�lߌ_~�J����I��c�c(�gI��;K�����]&�&}�ҩ�ҽEF�����typn!V["�1�,��0n�V���������f\H_b0X.� h�)�{�WNpFa������U�,��-O�}�!��QH/��d붔36�X�}�^�mVY����=>��f�<O��
~¬����H�++�B�2,�Q�"��j)���)Q�*�F{���Ē�f����g��a��8d�ԣ��V�����N�/*�s�6��B���v->G����R�G'f>mpn��Ծ\PN9��h�!?
�L�w4̌��9G.k �Y^ y��J�k�L�<Z'H������\�s9Ӫ�#��2$6j��=q� :8B-�"̍�� ��T�����o�l�4�e{�T���w��
�~r�=¡�fJ���.���m
�l�O�o�.���ԁ��#	�Ke�eXQg��Lyr��(-��u��8*j47|�i�eP�F�5I�����a�R�!U����~�B���ԽD��Ċԃ�MS�rϛ j�'�4�J���Y����%�gTSw���1�r��֡�6Qw�-@� 0���V�G'gm.- �����W�Z�����T���_�43�#�>����.l��!���BC;׮�=��w�xS��G�}xs��vqH�@�l�>����������^�� x)s/-l�ʭ�z�l"��	����v9�D��y��_A�CMJ��(鶬�#B���5׃�Dn��[jB�J�&�+�M/w��!mRl֣k�1�m�vE���[�M&�0W�����5���5��@���.�a F>px	��2Û8�x,$ʽR.���a�a˰ٳ�W?�I�Z��O�J�"���8��Dve���~3�+:���++z��3�ip�J�	�_���?�)���l�P#���+F�\�+�:��%<��k�ft�-��z�Q�w��_T��W�I���e9����&	�u��c����I�tT���'�Vu@�B���-�0�{�W�V��A�g"����<�w��K��y��fX���х=��֧[TN����)5�\��ߞ"䍌� ����-���V�坚=(����ޣ��Ԙc�h��u���:*ԃk�CM�5��:�2t�8{Ґs���rِ���|սgC�&7T�����pu��>t�>/����߂)!��	p����T���. ���+��g@������Ҕ�y��÷W��8�}�^��X���sG�[/�� �]/ء��.'��O�͙� ���O:��H���6��a!�#����� �)��M,��	1��$'�+�by��Q�a�L�+b=���e���:Z��f_��B�,H=��#sB�W�Q|�GN|�� �I���c�4d���j$���o�3X��-�K6����.�WC� ���9fHSG�J0S��2u
xX)��`	8��Y�υ�/�� s�d�\wZq���ZB���҇�!���C�Fh�}�EU�;���hR��.�fc,a��Y�l���m�� 7�ѽ"����Y�����u4�������{��(d�|Q�l�T��G�4�xթ�%.�$2��
�ʏ�yR۟�6�w��MI��8!��规�4��mk��*?Gc!��{	ݎ�"��� �ϙ�=�;9�'}D�lMT�����v�����n^D�z�v���6����P!|��1�S0֫�br�6�N��4abI��f��L���_]\��<b�֬��wvI~� ��@�N�oP��N�i���k\��&�4T�r��c8C�b���W/Z�krǁ��*6ع��t���{d�	!��1>v��:�@�c�-@	�s����?��Ͳ�!�5�Q�N� }�8h���m�����%�ı���R�[z`�{c*�����叛���@=�` �5�Q0���Lޥ�▀"!	�j"���PC��~�$��Z�)��f_	��L�i�e�̐Z�z^,*����+���yiI�(n Y�)R�K�.f۱2���!��J��m�����1�{��,Q@�9�'.��m��}�N]�լӪ���e�G���P8�4�+� JV#?������	�
�vJ\6�