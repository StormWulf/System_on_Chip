XlxV64EB    fa00    2f30?Ƣgc'��A*���p�����yfX:,���C=�anM&|�"���wl�Q���Q|���� �VwF�/�;�4�W�;�f1�58K�3Ɇ���-�� |�E�tx�2�!�b#u?8R7(��#�����v��ĝ�����禴�L�ԍ�v�xj�X��,�ʢ�Kg��M ����'#S����\�B�����y��t`�llDU|&���kإ�����p���l#�ڰ\]���U��鹪i0?A�bㆣ<�⑴N�,�dhXub�c��w��+.��v۹��5Q�L+*_( ��_�a����E�\���)���ɜ^
�����F��ȅ6nGXp����'���D��N���r1�H���2F�������b�񩤮䳖 ��"�J�nx�B�j��A\�]�3��ӆsR��AȌf���ya����cUC�(�#g��	k�pQ�tD�۪h�s �}�NYE��7����0g�p�u|��k��+Ϲd�8��4�����)n�B����'��4	�8߱�+��v�n�.�ѿpdf��o��Q�5��G��{鑵b��M0H؇mG:�X,��ő������a��J�S�Vŀ�B00oD���,�<�6���B�7�ǃg�e6Ə0⯶k�&�5̜g1�Y���V�Op�*�nN�����s��PλgR�H�H��4�ɗ?�:
�ЕdhQQ� .t��!p g�u8�hN��د+:�����3��9��DZ-���C�{��a�,�"��{L�v�ަ�x��r�����åa>�DyQC �({�|�6-�_���.dI`�)��v\(�] /Z�������.t��ǜ�&y`�Tk�?<;5��ᗺ9�1�=B�>G��?��B�����M�d�lA�8���QPt+E:b��:l9�%�Ĭ����y�:��}z���R���7U�LD&`jg�ֶyN��@}�X	ܡ��5��:��+���_e��ũ��u���"w����=�ЍX�T+#s6HN�]щm����.};����%ǌ${�TL��p���߮��h��`[�=�].�i!��,�La�b�Y 1��1���sħOFT
�Z��a�@s��AE0�j�$2l�!̥�O.l��].�V�( ����	]�15�,��.������u�YA e3����@l�B��A��<ݙ���9��L�vkrm�%1�[1䴣���:jٸڃ��P�}����Fh�����,}�К �Ͳ	U7?�����د��a���c�~�#��n�����U��
�:Yi��	�"�tl�X&i�c���˦��V�u>�Jgq
��a�����X�w�T��rȲ�G�^}KW��A<B��l���:��ą���^�h���3��k�"��%�D��F�F�~=���~JZ�C��E&�3-Dȵ��\Mһ��^[\g2s������i�i�/8��JI/�ob]-�����wCl���$Ts*Le���v�/���p����W�T�8Ӻ��H�g�]�W�m�b,5�v�x~�������$D�c!ԣ�]��?�wR�`q�q��.��Ai}v�v�s��^��01��Y�z�a/����W/X����Ys!kS�5�'�K���hA�t�vrнL�#Ϗd7�g.鞆��F?ˆ��=�C@�f� !ݼ4;T$���
A�����O�.!�r� ���>�+QR��^t�3D� ՛��ɠ��J;dv��LI�˅�-�j'��d��ğ)�u��f���7���|�g� �(p���Z����Ԙ��C���.1&X��2Up����4͌%�?;������)�&���AW;&:n�_��\08��ν�y�_�-���u�SQ���z���Y���\��N�0m�`j[d����}�Q\Ӱ�X�M�P�(��������GI����E(И��C�T�=�[\��&ܰ�����*���&��u����p�[8��g!!ѽ�7�sZ�J�KĠ	�)f�qìƥ�檰�䅿�i>��3#uJ�����!��*P�\P�AJ=���*� u�U'�3���<�0֛N�U�^��.����QO�Uk~<g���tEH����v�j�g�۪,��|>=BEQw*p����[�"|���W�����H���^a��F8�[..�ޟ$�����ۺ�c^�V���%�}���z�9�����=͏����Fjn-����*��Ƅ����C���Λ�{�Ӏ�&���3�?����$d��豟����,ݒ;���ĐڵUϩdc,���t(�b����nSzٱН~�H�E1�Ŧ����Z��0A�qru���nՆ/� �ο��9��;����M��䣼�ǅ����;����|5j��n4�^�X'�ٞP��E�{�iy��pA'_]���-ji�є��<�V�OV,���oT����a�.cT��� �k�ɶ~��~���N{�v�M��R��}wH�W\�(�S���fi�
�:�\ꕗF�pV:�s�ƕ�.f0q�f������-s*�S��:��~W���Я��E���L�另�sB~��s����6.|�}#�q�����1:Uߜ����:V�X7SqFe�����s��WM!5�ResmS����2��Ld
��!K%K��eV�|�(�)��n?��& �t�lk���)<�Om�`�����뾙��X=+���[Lx�p���H`^2�V=��j
�G�F���9�c�~E��*2�J���� {��]�A������C��I��"��f���[g=���N@b��%8��#��^��N��qz��҇"�"��L��#��V�I��OT(q�՘b����^s����[q�dm�'��Y���?=g�
b�Kw�H����H�h�~�FQ3��8f4�_�N���77�D��:1f�����`���re>���I�
�$��;� �F^�1(��Ȉ!��l�������IQm��A�B��6�Qj��8�9@4���O�E�tw�*MӶ���C>�㦖] ��C8�!���©cx�Ar�]E�bm͚�� ��G��h�ú���Kk�@H��tk�#���ZU�v_����W����@������&���������`���7������?�i��ZUL��GNHD j�f��X��\-*(>xK!-����rX���C�6ƴ�������}�W���SN�.D�[8��	P��G'b0������&y%<�(+�'�l����c��c����'�` kMu%�w4W�{��6\�/I\��5͈�@��..&�/������I�c�%�xu�T�Ýb���ʖ[�˂$��=�ZG�`�>J7&;v_x��Ṣs�:�Rڝ���8{Ѐ�ҾPaJ˃X��` �g����r���y|-��,����.n��ŊfdA����:n�ݑ��0dwQ���H'�ݍ�c�(�pK��S�-C����#1 �P�G� �H��2��	�p(�Dw��C�����>xƱ4�O�+÷Ǹ�������klがOh��E�o� ���b��MR�ad��3#4���nut�ϝ	�����`�h�Bz�������m�e7�ҷϠ�E^F�[9Y��p�?%5A�E Kd�pK ����44(8�K67��	.-c�é��k���j��\s2�J�)��������2b�g���߽�I9s��u?�+�#�K�U���Q]6�훢i��	�P�*5���1v�[JǿB��<x;��=+RF�-	�Y�+�kV��?��+n�~�p�霖�;G�����ѽ�%��EK�0Q[�����؋��/�*�i~�3�^����Jm"�^v�F��)�
�ç|���^�|!�o�2}*�~A�:�kZؾ�-�����#�I7t�A�lB9��_c����\�)O˗T�w��pX&zU�d�,�P�� 'A�r�R�թ�w<6�y��y3@R��n��ɍ=�P(|l�i/�n�:x��1Ǽ�)�p*���*t�kո���+MQ^�ޡJ,6���]t���鰫�������>?F��e�zp8-�4��1�v���/*\4���"�!~�K@ 5�|S�y��N�=Բl@`[1Ra��J��w��yI�w����#��N��:
h�`�������#�6���N'@3V��$.=�߉�)��i�7:x�ޜ\���b��|���#�)#�[M9�HF#T ��*Fyv��Th�y�gW=s:��8Jlz���eOxKM�R7��C�'���ϝ��$#���g@�T�0����5}�����6Z�
P�롰un��9Yl�I�ɼC�	g1��@-���"֑�>G�-����c���A���f0�Է��3`s���@*�Տ�4�ck녯��4��t����S���W]��Of�k����f�3��(!�0F�8�8k�V�-������:��d�g�:8]�,>�S,.�a��-���ϟ�ӡ2֍�0lP���֣f��TfV ͊��F@1��V��ԅL�4 `����19+�plf��z`5z����6��i%����YE�3�Ο�����t�"jy(�f�l)"��g:u�R�g̻��i�� &D���g�"�R�S�NB�:!UGCSf����O�@4�E��i�o��ʤ'����\w���m%���̴�rA�� ���D�u=��u��)g8Y .�9`��-=��Ҫ�n�gxy��7%��|6gk�Vv(Ls�ZR1��K 
��>t��"��b�~o��VrǦ'��%\�w	󁏈��X�^�bz<��d�|nm�Z`A!n�:���=$ 6iU-d��l�2�������i,�k��H��/#Ы�9^3ذ�L��Ռ�nnN�Ȼh9"�E�����K�(S��n����տ��?�/�<�J8%̹8GbN����?1�M�ߕh�Йn�6�ǵ;�����'�Y�S�N�7��5�	vX�Os�^y��TUt��ր�g��5���S�X�v[ɵ�,ڂ��Nt��.T�m����[ �gl��\-�h����Jڛu(�t3@�Â����D7`	�>N�{͠�!m�c��C�\������<���V�q�"�>b��A��_@�6�~�xL������T�b�\C)��x��c�]��;H��n8Yn톥^ K�-~Ϲ��Z�I~oGx
4�����������p���{�q�H�Ÿ.Z���K
1�P�����F���Tj���#q)��.� �pV�Ɗ7����H������Qr��'��u.�ȴ��ǐ����xBj��%�gҿJ3;PO[�Ď��b#�[�;x��M3�.�M**�r�'`��A2Ap��TӌX3i7j���(-Cp4� Kʢ�D_xLx0�Ҽ$�l����R��"�Jی��L�M�@^Eh��>�����hk0�)cl�b�wX���(�c!'烅rGmf?�k`�lA>_�p8�ꙛ�d?���{T��YLq43R�E��5��Z.�׬`d��ar{��y���=����?*��)���a��c���.\�iK烂���ml��V� @h=�Jz����^v콅;�����Oӗ]�82�C{ٙ�&T�r����:�[�X d]��%�7ͬ,�X�P� �t����{�43І���Q�Jp}9Ic�=��9����8i�&�a}5Ղ����5P�kOB�D��K�-��.���ԋj#��1W�]��wQ�x��Ȁ$��!��gS��;���DO��ч[���*K>�t���{���7:�U��<Dď:{�󽌫m�@i�C���q1[��R�ͬEp��ñG�6"��!(��ϟ�:��?�'�Z%as��=��?���?�2�go
P����Ŵ$KC�~�/?��C�K��ϟ�	� � ���x��_x`q&�y
���8�s����s���qoN̔6�x��;|��CC{���:P��ԁ�Q���;�n���g��x��%��D�Z��a{�Dm��!��L!X�,���mњԥ�!�^z���
5�c��c�S��%�'�oY:�O }7�:Xk��vw���޳5�����$�J��L�>���oK��*�ߔ\�C�F�ӟ��g<�����'K�����ً��.\�+֒-���,f�¥9X�p�@Ǵ*o�4�2c��f�g��JQ�3"x0Mۅ?Ϲ�NS1"����#��`�Oe?�N��f�����ނM���6~w!Z:�N2	/S�bf�组1�~�xT��lj�TA�����$��|V��2`_޿S�"�.Kˀ��P���s��GP&�8�Q��$�2&Po�!��?R��Ws6�	V�ֹp�$�so�D�x>��`(^OŲk$�-P��H�s&ƿ�H��rX뭙����R��F@Rx��`_�z��ZF��╩
LC�W����'�녬Ok����*�����$�Ө�d�[��H�@�n�iFnͩ���c}/8UI��Sq&�B$�ӏ�7������0��Z���kg�sٲR���}�xuY��d��1�6l���L��'S�ZC�:>�����g�LI�!.f��?�n`K����P�5T�� �^k6�$_f����(ގCv�C����bjD���W������č�į��_�)o���v�dA�*���`�d��/ʙ��
Q�tF��=�ڪA*�Z�}
��b���H5�Ǻᦍ�&���by�5sߥ,�h"׺�B9:�Fv��!I*zh���dp���y�>,�H��~P�'�B�q�<�c�hyh��߿ن��s�J+L]j�z�&��?�Q�Hܻ��\���wbT���i`���$��k��oC�Q��Wx����!8�#���̜a_��bo�� �7��n�tYv��sM��/���Jo#���PDn0{Kd�Pk]#2�`͓����cv7_	ͺ�\���0gU�Ύq�ٺ�^��R���Tg�!���O<B�QV$0œ	��h	�y��wtp	�5ͤ5�2&��ׯ�'-nM#�����[���2.ϳ�f�.�D��̮�$o�򮒁��W�!�o�˥t���#q�AI�!�v�OPo!)1S(��pR]�6��jl�yv~Y�w�Lf��H�Zs����N�w3l�)�go1��hJ��]���)w~�Uf����I�����L0@sӒ@���J$3�;�E9dL{?�~sՓs�3��iQ��X��v�Od��b�0yrt�J�Y.w�>W��`�_��yF=?��oA��؋�jM<�D=��BNd��̵{I| �0&<R?늅֤��sc~j���녡�v��`�Q�w�v�g�߰��iM���@Z��Z���'�)��C��ۺx�=>+�9޹O�N�"�xF�9ʹK $ ���	�=���v}h�f,���h�7;�'*�q���z�W��M�,�{G˰ҿa�
WL��To�C_e��7�'>�/�f��@S_e������7��R˹3�	jF(9��̀��j6�!Vg��I����@��|���7�EP�C�W�.��x	|{G�O����4�ǚ�ژ�^���|��)�	�k8�ꚉP
6���}�{��j����,�d���cݯ�>A��1L�떜��������L֣y0���ʿ(ݬ�qq9����?�wb����q�N��S�t��UleH�*e�j�E_s]�X�P��?t�#q��X�2{�D��:��R�?�Y�A����������L8c=N&9�6�S��_~._�uyvC��edT�
T
����cP����	=<���N��!��[���a[��i�w��m����7d%���@���ݠ1LU��S�귘t���h��B��|�2
�x|��m�4WMJ�����,�5I	�c���#Pll<A9�{!%p�"ȀSΈ��\{d�����(���&V)^l��������<����t�YP�T��O#�qLl���a#�?Y�`��	Nwi�:�t9�!^:t{�4c�����N����)�!0 �=6�̓��U��=K�p�����=�1l�G�n�psz�Cʾ��'w��8�vEHg9&l���ʏ����p�m�i��,k���\�{�}�D�o?��?�� �ᕽ��
�t"u��zIs/-m�L�"���Ȱ�x4�Zbi X ��:4����ZY>䄟��n����r@F��}��q�6A���Ǝ��u����k���G���>�pd�5��7m��NS� �K���g8�,AnӉ+9��o�M�ߕv9���D`a�y�(;;�*���8�2 q�!AE���r܄eP�V��қ��� z���H�8�p>knh���M�0(8�)�'r�׊�_�I@��Y���n#C��}@U�]�ACį��ﾵ���fD�֡n�n�#����jI�T�AOo��RL�<>�"
	�XU9�~�E�=vpؓOw����W}��*�����������בּC�Q{#����L)�R������Ih�XgJ<��đ\,����&��[�њ�L��>,���|N�q���v���b M��t!��&o^̧� �R��r������8�6�!�."AfЭ5��5��+'6�D`���#r���=�j\N�#��7���S��o��3e2@��u1�� �tVq �>Z�Kr{�ڰ�{�\�Ρ|,�L�n(bHf��.fL����D�� \)���خ�v�f�{?[wΰ_���yF������W��CB͸Dc1cձ�vzi��
)�7�_W�[�Y��7�4�]J���HL���L�lR=��xdl��]}e
�R�3�]7�
\�U40���T�sNm@fq�8�%/��'t�q=�f3�M�~�R����z�5 ��ᄝQQ��
bl�t�ks�'�t�һ�.7�[�C����\� '�����;�^y��Fd�Є�)N��.�����!�\��,I��I���@�� �`����=���t���{� �4�b��:��ԝ�>�����d���>e�yb��+p!�9;������z|C�e�� �ɍ	{��bT�;Oc��BFG�DK:�ZK�
�b�C�C�dA̗Ti�3�����-'��ߩ��1�-�M/t��>=M�=��H�qk��6݉����`�~e�8��(g輊SZ�̇���։B\�r����1_�h�j���%5/9�����@KXyשau���Q���?ʽ��7��n�F�z�����D���q�9���AlU����g!8m8���w���K�7w��\W�mx���6���!�ZA�p.�v��*��G� `�E���Bcmsر�fI�b|�>Sp�|;����a���nQ�!1q���z�y�|&+�F�?���I�U)�A6p�w�rw�c�y=;G2�&��	2��*l_ip���p�c���Qz�&(8��|l{�F����𑉨sJ��������Ι<�k�G�~݅{T���Q�4���6�q��)K_ҥ���g�v{�����_���Vx#��j����8��TWB7�z�����G�_�McFap�W�X6���Q4�~��7G�~>s����-���(�J�;����(u_�;]�B��O%��xV��7/�_��PĆ�jq �sF3�-�!�=��Ü���z�2���;��1�}M�\oR��{�@5i�/�%����;?��s�:�U"��������QD�g�����~���B�0[�:��V���e���\���*�2��{2D�p���u�@��\�6+�k�:����^�g&����ZrS�e1�Q081F-���G$-s"�����,�L�A�!Hw1���j��J_	݂�<3���(W�#u�"�!�x@w�T��E)��&+����ܐ�c�;Q�&�ɤ#U�-����V'[^�Jb��n�솅,���t�+��T�0��x����2��H�ۜ%&�Q�u�>�+�;(zy���/���������84��=�g��[v�3��,������I���~?�˅gra�J"S�b�l�9��jP2X� ę �.7��3O)��P|n��*�Ź�K�@H�7��R8���xN�3�!�YR�a�֕�Z-xˠ1KEo]F�	�|mv����W��A'� ���i��)�K� B�ɗ*5��r�&��`-�fHK�f"�^�����#����YR��(�����,E[���0�9�h����t�"gk�rTa���<8���V���Ul��@o#�����jy�_U���S����e��(�S[_[���J�!�m	�`��_-��Q�� :���?�7��f!2-�g)v�F֝�̃x��^l,/L/|�ML?�Q	�Iʁ0��Ӵ�n�̫���]~@�0��$oI��G -���,�n�� 79�IMn'b���B�?�\�5��<�|>��{�h�P@�W<�E���A@�g��6t�W��c�p�@�:?)���P���S�?��ߡ L��z����s�IS�	�HsiQ(�Z�4�d�|.�(x��Ks�D��l!�gy ���E"���Kb�/@qy|��b��N��+�<��=�~Hʔͤ�,qy�}D M��[lԕ��eS�^�1}�ӿ��9V9�.8π���ġ��?�2�k7R�al�f�Q�b����B�z�קE�)���j�oI�T�L<;[�����ՒW�2t�kh��'G�����v��)Z�>�Ɉ� _ף�9"�˗H���i�=�-�Vz�������jD��D��֢����q ����Aͭ>mz��y@����_mfl�1d;��ϋ2��y�h׋����*Q�]oi~�i7��&"^�v�!F���Mаhp�^�4r�$���R�9A�s"2��du���m�Q���!��^cDl����!��,ڼaڤ!`��#�O5�d� U"�Ix���
~#]�C.L��R,���4����q�gʃѢ>S���Q�k$����N;e��0� /oG��"��Բ(���ӟ?"W��i�� ~O���]	eoȻ�i4�_˲r���w�vj�A�]���
xi��d���6�q@4)9ȍt�=��'�c�=�{+DBn�����.Z��v;q����c3����1mm<ζ��y.0�|+O_�����r����V�I��:��m�4��`C�Ƃ�q�~��a	vJ���@ω����3_g�xB߬��#N>��:X�"��ws\�|�'˩˻r�|���]�݁`���A���:�yŲ'���N�&�?�%�/˧T��)��x>м�����b5h�P��5�V���0Ֆ�t���8%ZyʤX��� ��B����Wv�"y��p��~����62q���2_�#��{������P��Ze�R{5�T�]�3�����VN,�Ckub��b���_�1�xy�mڢ^�(�v�)�~v��_��Dl8A}�w��K�4`N��/<�ll��Ek˼U��ݹ�g��/�鍭A���_��*�}�z�h=��,�%JwSݳ.K_��k�2�e���KO֍� k*��
1���o����D�`'}�V�񛸥T5P_4P��~&5�֣��X�֞}�%̪J��֒�i�f��s!�y�j��ҋ�nA &R%�ui!G*�h]��5�YR�w.�y��2�
#�ܗ��cd�uWC�v3f�����J�,�ow�am//'��g
z��������Zö�n�(��FpT���z��.�f��L
�����s;,�4�XF���,�dK�刓s�����Ǣ��?�!�q�<�~��oɴOF]@l9sb��� -��-���|���C��~f̈�k�|ns���I<;�&�<j�{�G+��!z$qz�S�ߛ#;����9�`78M\�x!y�lP�=*0`�n�9�2�,%kYn�ZO�޷LiȐi)��)y�t��-��t�w���'P�*��XlxV64EB    a4cf    1bc0?eu�
�m`4��<�`)g�e`+x�t��޲o-���1�����wc�bշ0tss򒖜�t���#O�8�>��*��Z�f�M�O���<z���̧w�
��q�E���xQO�iʪ�AhuJ��}�/��N�,�L��!(+֬�N4y� 1��gŐ>��Pp�7�_��GhS�mH_������r�0`�
���-���a�.����3µD�(UvN5���Ak�r�
�ڷ��n�>��ݮ<}�sn�$�u�l���k�2�m��],A�k
�B���+iq�ә��5}�J��4s)���v㇜�V�fzP4�~X�K�<ڦ!Z1�"�~0�*���1�<�O?�-)ׅ|.�}!s��XI��?�
gl�!F�.�XC ���h"*Ԟ?�E�+W�����1ԯ�-���$�U��eHw\�ޗ����������@-d\���yx���i�l�k>���kW���p I6���A�}���G���;#��3Lq$��p�	�"�4�Jc�QU$��M� r�-y]�P]����\�[���׬Q|b�a����[:>F��>����t~�2�ϗ�Y�NtS��v9��������)<������7��*s"��"�]m*����L�s��v�E7�|�U����q4l�@O	�?#���
������De_M��s��{��8�M���˛�#���SB�=�GT��7� ��`ې-��<G�u}�f뗚	߇hPv63�=�:���MM� X%R��65s��N��ß�����m)c�j��Eq�㣷^bV�}�u���*�i��m��)����Db���i.��@����WG�����s�jË'��OmNlF�*�io1��V�vȊ��>��6s+mܘ���q��S�n���2 lDP>\�������7pD2M:m-�+��a��)C��:w��a2��TS"��$�C��V�E��:��d +CU$%ɶ*�7�[�48�^7�-�2s4_��E�G�9�L��QF]RP�8��&jZ��˩��VU��r��һA�=0MD���� �^X�1��k��$�إ�k�Y2<����w��܀��Y� =N��c0a��.�7�!�0�K�Q
�?�a7�:�jj��1��
�h��YM�����J�&����{v�>淫���ql *hOe�u�$K.�; �.���5]�C���ki�6a�-�ǯ�m��*�p��H'%�{���K(���Ł��f�p���d��I�C�ѽgu�8���J����|�Q렆�u��oz 8�^[�0���(7]HFC�G^�N���+J����74ب��[Z�'Ԥ�0��\�������}P�jbM��`m4@e�f��#��&�+��#г��:2��2��1s�3���n���3��&����s��ddR�8������5;]�]��/a�$��5����Z� q�S�P��*&�*�T�DϞ(�R����BM�}����il����oE��]~c5�)!�V�����]��P�k11P%�(��0�?���(ᵭ����. =:E�@�g8v�`�%��zTܚf�p'NA�@3�A,d�-[/��dDV����B��g,���HhĲ&�wuN�)�N;�I��a��~l�ђ-{�s��4�h��4sI��h�-2:	H��U:!��^����-�f5��/�+�`�X��o� à�"c��\�&	�Y��5!<�z���Dc��Ŏ<O�S�o�Ѓ��N���|2���͍�ET�ѵ�%[�׋��#�RJ����P�ڲ��׈a�����
���W�CTm�a>mH�K���n��������R,�$�lE�A"%~8�W�XC@���<(�|�`!�t
I�B���z]0��s��8+(\�A�ETrY���K���1ޑc� ڭI%�2XY����	���.)$%��A�M�j'��1fB��Kc+\Aj�S�c+�V�K��#�##��'��FK��K���nNƴ}�*�R);/�(�pR�rnb�>S�X��Adn�!�0�,rWm"u��%�m� ����3Z�Np.&TH5��R|!�|�O�z�"�)I�+ڍ��mvg3q�x��8�]��K9B�-�r����>����:t�ee�s�Λ��1��[Cz�q/kH�q�{�%�%�����^
�o4J%�T�>xLI�,���8��y�^)D�%�;�޸�Ɔ�~��M���#��,W�ȵ��6�[��B�d�>k�d����]��ǈ�<o�xVR��m�%�+���I��|���;KY�[1���j0�w �O����G��r��+r��V%����.u�v�-�r��]���4�MI��ǒ:��_I?�Lj�hx_�]�P�׎�7����j�;�~��E��C��ҕ�읥�,ӆ�&G0�v✋���$3P2p;��otՎ��]|g�@�o�%��og0H�R�яҋ�g�|s��w���5��-K[��&����6e,!0.lx?+D��� i_l�jR��E`X��M�����Zow��Y���~�Ϙ2m�{R'!����n����ֽ`��
�v~BAl�� ��&�2��8�?ñ��Ɓ�|�\m�6�oGZ�G�v�{ϕL��]�<L��RB(����"�K��pf�x�|�^,�5���'ث^����栤Y��p����XJ<�PT~"��ap���&� k����M�����s��^�Xc��8�r���_W����j�j�f�� 9h0Q�H�}��-�� �ϫe-wED�Q���,�A����EJ w���.���^m��S7�5���'Wau���Q��r�~���)a\m4��D���mx�9��8=2x���vp$�]p:�m/����l�73�{�1�:����
i6$�)4X�r�H5�����!�v�]J�m{O��**�O�i<���3*o���$�+J�	�j��O,O�M�e��Ro|�g����F�C�6���>���s��K�`h�a�����Z��?hm�l���*��iA�0��>-:����AՋ�-�-�L4�y��R�c�8�e{i�<���N!��@0�H�V�*y�kV˙�vQ(yb~N��AW\m�⏒��|+J�8�}����%�W���֥M4�o���y��>��тʬ�r B޼ڳ�ǸY��q=�( $��¨�S/�����g�����,�0�R*��ڹ�E:5���WA���H�#���I5}?OvML�V|_7��9^��s�Y\*��C�G�X8HN��pi�sͺ�J�4!�v��Ņ�]δ>�ĲF5�v�����<Y\��c������cf[��O4c��I�A���y-[x3��I�1Or�)�tg �y]A��.�&���	�%�!�U�=igV�-��G]�K�MZm{�i���..�K�\�!�ԕ���D`<&�0h$eI����R�F���9��DO�_�w;\l&� �0Xc�c6J��s2��
f�	.F����dԊ��ǃ�����4u�3�	�����D��6�J��Ih�4|�Q�~��A�Mr��7~��&$��#�l�`v2ה2��!N%;��Oy�GP�Kg�(�,�39��
�9�gk��i�P
9$Ɋ��I�i'���x/o��>z�D���,3QȎ$�p�5����7e�R�ee2��I�cə��c?��ye:��K��%m�w�]�!Y�[zl�':�qY���kV��#�a����o�U�#ǀ�I��6b� 榴�&dv�i����3f��~���QC8�q�f�X����i���Z$䮣M#&�,�?f��Bvo0�+	Mn
�5(�k�w�F&�Y4��2	*%��r�ԁ�K����s��H�Y��@ 3���/�,|YH8��T�j��Hظ�������#�fH:���K��� ���A���1L����8�?���b��^����@��O��᝻&
��IQ��c#�Πω�u��/l�լ��=��ɩ��Ӵ�slF��|�����̧���X	D�&!V��}���[�[�a��_�Vh��4P`��Ղ�z~�Z��Rp�@�Rb�V;X��rҖ>)l\e�0��\��������]��& ��i��({[�b�f���:���A�i���iEZ��ҝ��E�J+��ڋ�V
S�7�p���^�'h�+�*h�u.aS�����9�I܏14g����/���O�뾗k�ӄ��}�i�@�U����Ү�4�>�.]��Or����O�&c%�`�mx~t�e���ŏ���l��L�USv��&�"Mǳ�?�ʴ�P�()�O�e��MKH�� ��{�ޙZ<mg��3��C�ЅD��6���/�K#�]$��k=�i�s7-Ί;1�kw���:GqMG͐��D�d�B\.o��,˩�W%�%���-�REH��"���J�j��[�iy@�L��Gr���t9F-��)7��u܎rc�~�본}b�1n������nVJ�L�g04]d�Q�,B����ǳy���`@��8a�[Z�y�����T���Aكk=��&B�4)���dJ�� ���G��$	gLxF��S�����$s[ �e�=�HF�����2Kv����8r,�~:��O �S:�HB<�o���{�/��.�r���`]�O$��O��S���ō{�ȡN�+~��R�o�\�Y�f���J&|{�o���m��]�18o����|}>�gk��X���_3J���<�!��EY���e#]�J�Y���E�` �#�#x!���b[�;���~�Od�zԭ	)�+�)\�B�@h��Kp������E^=��~�
F�k;No�=$���g�V³��Qc.�yct~�1`�W����|��0��sT���*"���REۆ$=�v՗+M+x�i����-�c���Y�kH�~��$H�����O��8�}{?�x�-ķ[�3p�B�h)�<+Ӈ;����C�b��+0Շ&�>/�ߡ�XX�	<��@���)ƫǜ�}���G5j|�}+9��0��>�5ʂ�'��|J���5��3HH�ޛϝ��Q�7������S�6Fǆ�]��d=��Z�H\k��$�5��1|jd8U�ߔj[� ;���g��I�Hȯ1��KNJ�2|�F�j[�yى�vc����Ím�bD&?�TH ��4�|2� ו-����l�G4y�^X�b�����b�,�v�$�C�@��ݯ�ތt�k1$������<�1�ť�3s��K��C��@��W�V�)���
ig�m\�hIj���w9�B�>��+8�\�Ѡ%}��T�cKN�
h�*��O{�n�Tc�aQA�/<�I?��|�.��L_j�����6�]�o�Y����㾱0w@(� �g?�R�+=?�h2`*?R� |��I�+e�?J���X�f��F��ވ���<#e��q��4�2��#��jGf����3;�����3FEBXI����goX�ƫ>	��e�D��Q���{�ނ^�J�!~��#�q��F{6�7?㈃�0�7��	;ٟ���٩'�#��n�V�l�Oo�`��n��V�!�^��j8u���K ��n><5.$�����x]�l�,�5�N9Ys�ؾ��8���8G�A�����S�j�x �"?w�{�.=���FaThG]c}>�Lz���(~E���\8��W�p�R�g�E`��ߟ%�ܲ�FRNj��
V����s|E#�z�T�ba���E�>��5ȨA�������_����o(�Ӓ����=�q��{�?�.W^.
1A��N3~�J��� @%�q.�V<&8y'n�����'���
;�iK�?U��#������@C�A�@��q0JX�+-e~��Z��x;yտ��1�^�ȎՕ?E��Y��Y3~��o� ��z^f��Ն�!Z��N���B�l/�%a�o�������Dl/(�
F{ϥ��`t���5Vb<�����H4��2mM��+2�=�J	�h3mvA���>�Ӫ�H?�M v�kGdV�sZq*]��vT�ٓ.]/>��x��~+���ߧ�Fc6���z�LD# �T	���uݲY��p�~;(�b�n�Y�ֵ@������:&�������~��բz���ԩ�~��6�'�O!�/D��R���(%)�O]��(�1��^8�L�Gd�����#����~�ԷJw���X�'�7h�'�ϨBU�p#����R<����>��ګ�@���#��w*k�@��Vi���|u�G�3݋��&� ��Í�Q���AZ�ļY�/N�'n1�5O%o�a)���]I��[�jY�ś��ڡ���L��+RͶ����W���':����w��7�"=������f	"�a���<�Jp 5�b�Ղ�"�qюo!h	3���-�Es�x��!7]˻��s�>����$&��]�;Q��3�vǧ1F\���<�bL1:(�����m��BзG�M�wj/��y��~(Ȩ/����>������[���h�����gQ�A�씵���EX���Hk==@bu��l��=�P� W1�s��j0��+�ojq��t��5D���fſ�g�_K����qX�Ԩ��6[[���Q:��1q��b��%�&8���>�hNZh;6&Ƞ4�X�St��[\��O���nX.VIFOe'��S`��cw������L</k+1��1_Y^�n#*�~���k:\F&+�;(v|���� JwS���xT��M�5)�����ͩ:ex(�ֺş�<4d��>TjY{�������lsИ��o��B-GI��A�R��Q�UODo(,>e��~<���j��kw�	�D�e.3E��M�w4� hJ���^�C yR���z��%���ӯﾫH5���D�8��A�pyB�y���@3@L�ۊhK=��gku���In����9>���6p���� �4䧖<�	�� U��$�Bd�����D��0�b0U������"c�AEB���cv�N�bZˋRt�ɰ���n�xx���z��