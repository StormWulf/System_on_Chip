XlxV64EB    32be     d40��9�7}����@Yqc�g'G��fp�l��p���� �^f0�W׃���,.���v~���O�f�r���\�N��0"�ozDs����JwS�4�0�m�C �D�t����dtQ�:��r��+�ü���r�_�� vo�6h�OͳPIH��bi$P1�q�	1�_����LUf�Хo��ʴb�	�V�f�]}�ß�V*lG�V�՘X���,w�V�|�4�>�j����w�aB^1R�`��I�5�1�6��&�:�|��!��l(�\M
��sP><TY#.2U\P�k�т.�a�]Z�
��Y��:ѱp���Z%�F���6J�N�F��t�h�㯨��N�#��Vk�C�R	)?1K�SE4���ܗ��~
7�w�b����(�0$$����&��0_~�Y�IUY�n(�-[������%9��xZ���(T���T�,'���jWL�+���cb� =o
�w[��_�G�(n;b����Z,��6�PYq?��h��#a����ܧ��p�舸z�t,�ۚ�l���C��0$����/��ݼ�"L%2kI����=<6��»�%8H�B��@�Ͼ�zq��ob�By�H�+k�rP��_ᢊ'p�p�Zu�������Z�gGqgf�d�{1�f���� t#���98�����oo�6I�H{:
s�ṵ��˄tKT+��9+������f\�]�$�>��!*�'N����ӾՐ��02F���8��W~���`HQQf��7�!8y�c�#@kwr)2j����'.��*�4Z���77v���.U��w�����@b�Ry��5�Ҏ!ep�^�e%L�p@¦�/�����Rr��|��%A�. ��oB���\��	a��k�Ĺ��k)!pa��"��+4�r���+4@
�����(B� ��!���b�ͤ��%Da�{u�æ���F��3�L�l�B6�����U�r�qc&�[�HW4r�i
9{&�G*y�~2k+�v��7�߹C�e4c��@؀�=��X�/ڀ	�"з�qUka��/腒��ܦ�4
��{݉�&��U�2�d�+t� c�r�8ΝX�A�@WA�p���h�$I��:!ڡ�J��U���w����~j�z�q��)�`����b"LB��x�Jp�ؚd���9�z�܇�ɐ5ث���Y�i$/ȕ�{]�WiOq+�v$? ��6�tH�Ym<�5aK��<kw�;*���`;ؼ���h�o����B�IA8\�R=jϼ��nh l���,0  �����A{f�������>o��q=�����.����Fp'c��<$ �����*�]Us�B�>d�B�y֟��<����OJ��i�&Us�7;�zaO'b���f�&���k�=~r�o7a�6�Z�f3�,���L�F�f��� ��Ҳ(U@������o�jS�G��=�T9̭���[!�m�3N|�7�9�����x��R
J.��W������a��V����u똹^���D�m^~a��ĝ�+������+�:;�g`W9}���&7K'}5�8W������Y���>���>�S����ÕVo�Q�@�	,��#�~F��2��K0���)L;#��,�i�Ne��#���Y���ځ�Ziۍ��qo���^H�R��/��C+������Yc� �Ku���oX����1P\���<bw#O#P��r��7�F��y�1�+�(�K�s͕�n�B�H����
���EU����ݻ�Y�I��,鳂e; '9[*��)��X���A�\>%
O@���^�����=���$��j��x��Sdg"��jev�@�Ky�8fR�Et?֒6�U�;�3�נ�����"ci�Mf8e[T���*��(���&|0�P�4KV%#xp��,{�;*sT-��� �y순�ũ֣���e�E��
��ΰ`���{Š�\�@ ��{�Pr6���g��Ź��e�f�pc��v���k���]�d�X<�]X���UrzQN���4�W�0K4y����}1�\^��?�X4���ƪ����Ӽ�&,��t���{叠#����Z�f`��#����N�?�C�?nTuk$�eLXr�r��b�݋s&x�A#oTAn�'ˇ�+�ǔwK���xO��eu��<Ō2��'��A�n2q ��+�]��6?m��E`#�6|���B�6�,F��N�p���퉩{�OL��y��O�N �ޙ2��D.�7ޡ���q �8���`�Pn�떴�,�&g�4��R�}::J9ʨ�D�~2��G<5���� hr�5B��q1�qro�N ��)�o0i%��.����+�9-5[�W �h�Ύf�K1�u4�v���U���R�̗^�e��#
k���*�����o/6�K��-�@�J�^��]�-�f�,�ʼf!{�<y8,-l��ᘊ��~Ѥ��4s��j��"�Q�q�$����<1��yܿ�L{���g��ϝ��N)��֎����m���F��o*ViKe	ɧ����>&���X�
�E�i�Bmy�$������S9cE��N�v��TAر���Ư�;;�w���-�.��w@ӱ�
l���N�i6蓗k�`HP�:�~���-*I������yt����T�[��ϓ��9�����������>��4v���G��3r�_P^��(�a���c��� ��ѱ b�������l���e�k���FS����kk��^J�';���f�Ax#]��V OB���|�s��b�3�4U,PR�k�?jmQS�����K��8����Mūo�<ɤ ���9D�\PP��_)���I2Ѝa{���.^�~8cC�5��5��BX��K�N�ڂ�H
�- �]0#�&�-����o��Y	g<���+,0��y��N�خN��A��ѧ$�Ѱ�����P.%���zR�G�n�<*����ʡ�.�A��@҅ �^r�ȟ\��Ax3n�Ҕ&S:w���>��2 ����}v�:v�b�P��'�7���5��ep���K\T�����lf_
2�����8K� m4kL����Nk��ڧd$F�Ql��N�r~�;��Zck������"$�\����s����%�P��ԱB9l��{�e�[�������T��r�»>����ͤU_�{=?�LE�]���j��B��,� �.t������ܙCm�1w��=�CV�c௩��-1��oi���Q'�ux	�.9[���c{mo����;�*A�x)�F���Ck��$�na�S��n�F���R�kG9�hM�Of��/i�ڈ��1w�� �|�١����/��D@������3n$8�hN@����T�m�<�