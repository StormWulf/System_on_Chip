--file: proj2.vhd
--Authors: William Putnam, Jeff Falberg
--Last Updated: 9.16.2015

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity proj2 is
	Port ( reset : in  STD_LOGIC;
           clk : in  STD_LOGIC);
end proj2;

architecture Behavioral of proj2 is

	signal divsig: STD_LOGIC;
	signal sig: unsigned (23 downto 0);
	constant cblue : std_logic_vector(2 downto 0) := "100";
	constant cgreen : std_logic_vector(2 downto 0) := "010";
	constant cred: std_logic_vector(2 downto 0) := "100";
	constant ctrans: std_logic_vector(2 downto 0) := "000";
	type tile_map is array(0 to 1199) of std_logic_vector(2 downto 0);
	signal grid_map : tile_map := (cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans, cblue, cgreen, cred, ctrans);
	signal mapindex : std_logic_vector(9 downto 0);
	signal rgb: std_logic_vector(2 downto 0);
	begin

	--clock divider
	process(clk, divsig, sig)
		begin
		if (clk'event and clk = '1') then
			sig <= sig + 1;
		end if;
		divsig <= sig(5);
	end process;
	
	process(reset, divsig)
		begin
			--if (reset = '1') then grid_map : tile_map;
			--elsif(rising_edge(divsig)) then stateNow <= stateNext;
			--end if;
	end process;

	mapindex <= std_logic_vector((signed((pixel_x)) + signed((pixel_y)) * 40));
	rgb <= grid_map(conv_integer(mapindex));

end Behavioral;

