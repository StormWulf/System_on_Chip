XlxV64EB    4c5a    1470�/'�R��e0�K��Wy��7���;
ѳ/n���)��[�H ���^`GH�jl$9������{�_0�c��b!����#�T���2M�xhá�8�j�N��̝<�F���)J?�K�����vmM���3�ΝL{��-Sw�9�Z�"��Uz���R7�4Lr�%��ga7�o��i���K�O��Z�|Pw��i���1F����I�+%��k �s�H^��:����4`Us���]�,gl��a]4�r
.�"���pLY�Z6�҉~�~�f��Ha�ca{��,��!�C��$tc�����a�\�4���Ƞm�Y)V��*6-}(�+%��]���y�]��A@�SV����i}�nF>#3�]nݕ��4V�"��n�'��l>p���2��ʒU7q�����z�!��HI�����rB�G���� �"�x_��y=�_����X|�$����<�.��C����&vM��z�3��3�w�-�p栎����;jC�H�?S��A�8�?�q(������"sq�w
�/����-x���<.�1�^�Q����#֣A�8�ss�rsqP��aGo��q0ک1Z����|�+U������ܮ㝳/RzRg��|4�Ί#q�Gp�m�٫Ļ�yC����Z�~���N�TOA����ꅂ�1��3�B�Rk0W��w9P�~T[�s�q�4�s�mZ��P���T�7�>�q��h�(��t���xy �
]3L��/��D�:��@rd,|L0�e�KW�*f_�����5C�1����<>c'b��[FFH����ꦖ�Hj?�S�z�K"��[w]��T�>��߄TCļh��@��fJ�-c��Y����4r�:$������A��):����%�_ X� �'�g�H0*���4�;/�@�6�Q�S���Ǭ���'`�������w���2��>A��0��;�v{��_Ѵ i�Y愡�5�=f��� ]M<!e�c�K.��� O�+;/��c����Ʃ���OP�2���p~oZ�yN;���%����`<ua�E�]��N����/���i �G��VE�..�ΘL� ���t5 �QF�d�@��=~1?�J7�Xǿ�D��Em%��<�0Uvm1���Y��-���eҾ>�T����iݖ@�R;6*p�$�`h9I!\Tx��eT)&�_�0���M8l�}C��s�'u�����A�d"��-����h��e��?�-�D���jNLW؛��lh�t���[I]���żq�,Oq#��O��L�ׄ��6���Hk�8JY���hn9�b"� ��w�����qI�4Q��8P���S�`��s���"�[���V��%�� '�}�2�B:��"�6��ǖ��I0	!�b��A��?Jc!M���$�ٕ5p5� n'?�i&w{�74,\+⿩�'�I&<�FyRw}]�?��`wQၟI�T>�ٰI;0a
�`�'�G�鏢@启���3��w��kI�#��û+:N�QO����|��(*4�!>�(��	.a1J�p��9v˩�G\�x+�jh*+^�/�Jڽ9����ܐ�j�(���1x������:�P�]긣���^�!���1���Ū������{�Z ���q@��Kf�h�OeZ�%V�����/��+�J�[-�g5�����Lk���ҫ,߁�n��杴��6D�ص���V��/f}��%��������} ��g���gf��7�p_���pjJr���[\h#s�l���F8���Q��%s�Y��Ҝ|��f�m�
���ҧl�+�ܰJ4]�y0�XV��J�3!T[^FG��vd�T��;��� ݶ+'�\��V�7]�w�'������.�s#����D%�`4�ԏ�W�� a�/#@�5��W ��솹ah�|r�+�zy�[0���c��Y�a���b�)��F�$��ޝ��B�'R��iLt�%�׾����QޣP�+�O:�bI��|7�Ce�c�;�?#W:6�z�_�Y���U��'h�j%Xc���ʜ%�E�#��S�HC�h�?�<��[�	y5e^�σ"*���%�d+bJ�;�y8=��s����V{�`�/*�IހW �����'�h>yE��d���4z��]��lD��x����t��Ңk3����*�@��3��V� T[]V� `�D>���蒗�I�nbp�����A(� �D������q���B�ˊ�^gȝ<T�'�S��&��[���U��%H��TnQIFd��%�]7�cL-�����##��F�%'�e��$)�> )��RPD����Ĩ��/FR��� ���kO]#MI�Fyl�ɋC�u���� ϐ6}��ݵ���yX\
l�D&F�5��b��᯴R���G"')���\̪���N�Ðn�u�s� �ÙBً)>������hu�ύP�CzC�0V"�uΧY��<���h�A���	[�Lѿڼ?�miZ��ZI�z����7/���" 7{��2\v\�Xz�ü�Y%�E�S����no]�XsG9(��n�'���w�0"�7�H��3
Q�~�p��|�����\d�b\�,R� �Vl��FF��m�a� .���w+�w_/��l����G�@����~����,�:%�~�r~��^�4�_����j��[+i+��#+�K�L�q��rbK��=X�u�|VU��=���ޙ�����d)��&�*ϡ�4��	��H�E�"��4�7�;�E~�ڹ0�����1�ԎWó���>�������[�|W��9�-��%h�0��<�IT�Gu�N��q���������Ԓ�R��� 6Uql��d�vw���ۢ�!��0�z׏l��RK4B�9H@3�z�D��bٶi��c|6M�W�gmP*G����΁�J������|��TLR���0ax��ͺ��{=�y���Ό�H��Gb 5�k�FO���5��vL��шC��r�ʆ��<�&.�3�8��O��zl�O�9��s3���mzO��KE����W�y��|��Kͤ�v%R�i.kǥv��=��Z�6hv�e��2Է*���\S������J����<q@Ң�~��,��l�X�&t^����䫯�]���3V��N��hw��*l&RU�Kk{�L�V�5	�e�l�0V��+��n6�.;�V�11��7����U�]qu
���ޖ���m�v�!q@�,:�f����'�hT#C����I������4O*�6w=��!=�[\؟(�J��Q��K*��:d�K��k�'�^�ҝ?��l_���-�h9ͳ�1}��U2n�b���>9�on)(lqԎ2wЩ���n�ʼ���@U	D��s��ܛ�����ש���=�;`,�8z��ث���`R͇�<����KYQY�⣟6vJBڬ� ��.!��,�޿�1��=a�jm�������WsUo*C$NvK1�x<��1j�vWR2�eH�ji_��Q�����2��N8j+��G�89B(��̕_^`���ģ���e{�}��1 �^Q`����4e`�*7`'���P����8��K����g���7�*�|�
rY�l�9(#I`[���;�,�IaG)�鯧���x��z���M�f��<��:m[=��m������[��_܎<J����`rs>�lYM�M^<�TpҺ�O6�Ȇ��=}�v �}a|�ɡ���9�Ua��ᰴ���4{�u�S�o�W��){7'��[(�}oM�	�L��A]��W�΄�pFk�';����7Z��R��� 瘼�*?xβ�����֢.�"��s�m?�ukwE�U�����'C����|WQI7H[�KL�a�xj�����������q�K��˝����ۮ���ķ�ՙRH����Z�q�ZX�F��R&�@gQ!�W��G��N�ڍ��=�JE��0����y��|=W�-L���U�պcY�T�f.�Gi$*ڲ8SWX��]�[��LFb�X��-P�`q�l3���^_��J�@N����a���.���-�_P��PϷn+�N<q�V	=���+)v��Ճ�H�� >��[�\)�P��1:�@.�v{��>,d��������n�vC�n�g��چD��)�̡��l��#�)���8;�l�DǇ��]�}�>�;�E�#4�Y#A�(�?�b��跣(�5��N|G��(ȩv������G����H�W�eG=g�5�_6'#w�d��'?�V����&��w��+�r�ë�&Rm���}=a骓����D�7��^oL�����+�1:7 /a���'3��9~�j�gA���J��i�'�AF����3��Pw��a9Z�]Ꝺ`�̲E�+@P����~�WV|�
�I�������[��U���Y��k_`4
Q�6�W�urQ�nJ�&ئq�ȿD3/>��k_�4����x�ku�%W
�~>U�	C>UD.�j��sB��Q��iv�u&O������Q�rο���y'D%��A�^������� �QbN���@��}���؂��ri�Ys�H�F�ʦ�Ցa�ܷ�ֿX{���x)��p��6lXx��c��W|��y��KA�`u~e��!�\G/��Xc<v�b�a�؄�o=ɀ�(�hU�t�/�~>�6D��؀%s�(<��Z�O]��2٬��mWhbϢ�>�?fĈ��hJs��4��U�8�İ&��,|�@��b"�x��,��_�_�訧j6tV�E�$[�[����̪�=����F��W�a�1�TX����E8݅�HX���<�gU���Q����0?��@0/uP�s)pzPr�A����ݯ��O3��H��=nb��i�Q� �	B^�ةU��':``J���g�唕��Qp���t�hI�2�����n�W�.�n�9mNvy� G��Ÿ�$�z�׮.����u��x��0dO�pG�,�;b�ln���n����{3�.�r��n���3���V� �_�SV��R���pM�U����3?��؈��~0*d~7I���8.�޲Ղց�@?�v!�6��w�.�G�K��Cw��,PMA����������&�rM�/g}u�G3h(t����X�N4����`� c1h�G�w�0�{���R�_-^!e��u��Z�><p������-�ȓ��d��"����