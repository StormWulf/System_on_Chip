XlxV64EB    191e     9b0��/�4�&�|�ы���i��,i,i3�c���s3Č`|�AC~M�9�*�3��b%��'�<�
�xq�`�G!���<�Y��#F���.5�:��Js&~�z�EK(�k���1w�F��t�4	���<S�[�毙*�w'E�WRz�}��� �D��r/x3su�޹�Ղ�`�>�#���~�J�L��X�	'u��U��i�]>o"�%hbڠP�����eX��M3�@ˋ�^����&�W�HљA
I�0���m]��R�$�	������{��X4����!�Y�@fK����$�ߨ �H6|��G�̠BSsvƭ$�\�ۘO�ԪGoC��S����N(��w��j��_U_h(��f�Ɣ�S���p�����Pl�w���)/Ő� �`��k�(����;%�C�W<i�Q��ur�TNX�kdGX�f�����=9,��(�# ZO�p�J��g�L%[՚9Ji�jO��e���".6i�Zg��b.:��kS����FqOKa�.P���p?i>�������QI�(%�n��S4͓i�&G��e}�q�|�;4���4I<86��Dn݆/�1!�V�<�>��q���-�ʓ2�1��Y�ef�Y��<@"���x<n��Q�ș�Ñ0� �㭼o���^E@��H"# ���#8L�Kz%AΧ��3�,t����@�J�K�(�^�Vs�,��V�>�* �Մ�D�S���,"}��k������P����K.����c?A�y�v$��I��)�h~KT^ML�`�<9������3�9���~�u�`B�s�{�
�Y��� ����7%��}UO?�ػ#�2�f�0��r(�`)L����ҭt��L�Y��"��Fu��I�3����Ʋ��a�c�r�&hq5����!����0�O�	k�����RR7X�76�]��/���u)�ߦ�-�@jM%�AݙS�VoM�mb���8��4�tF�*�>z���,g�@�O�����}(4}��'ق�yl(˳�L.	�#�dߏ�#�h����>M��ܟ��e"�_�R�98!�h���R^t|��1��S	���o��U>S�̾q��k�Ъ� ��.ʵ�/ް�`�R7�{��/r��m��ſܟW@yk��X��a�� �Z�8j����>�����eZa�M��P>*d������� ���D�@�1A���g��k0(Yq&%�+�����˯{�h^؂d'�_�] �5(U�O�`����*�N��ke�d䦏�_{�'�v<�"9+�j�����ֆ��I�K�/Ro��Xw���A��:ի���-�эj�PBL��˪�]��s��0vn��Ĕ䢭��Fm�ѻ��$`5�x���L�˫p�s�q�dy���rϗ�e���	�:`�$Ĺ�m��ņU��c@YϻG�݈^|CY�Ml;���~�S ]�/և�SFYC�	>��P�gX�w_�RF��4z���S���Y%�sQ�_}ʋc�\g���H�����
���������n�	k�J%�z�!o}Z����d��ԷH�/*��X�!�"���� �,��g�m}m��m��IْCj�gZk$3�-�L��U�J����GF��46:\;�2���h��L�H�v`_����'<B���f�}v����鸽*�d](�O1(�	�ѿ��os˧=���n���_lv|��fg%0]%��ut��d����ÙP��!e���Z���u���)��"u���}��Z4�9F���[Yǰ�54i��~es�`mQ�w��ש�
��`U�6��Е�=��_4w�<9uY0f�>�Wi�������?h6�N���n�cI�M
��OB�d��Ce�n�L��*�!�*���BH��U�}޳��ê*��Y�S ������m� �(w��\��1�ɖ���YRV�{d10�zI ZG�N��d39)p�?��OCTg����6p�w:Y�����*�����%���p�=˼�W�qs���&+Xio ��{�ŰS���5:�[�t�jA��)�"@n��l��|��s��j�Xh�ۑ#Ԩw�6�ZV�D���ִ����}�l!D���'̇'�V�����%
D��ǵm�ʃ=�8	����Õ����۶j��Q1$��#����?���uȦ����<�l\�+֥vO�r�Ѭc!P+��������=�	WH�� �p�.O�	�A�p`(�gO��2� �H���ѣ����˫����7t��*CS������>�ؗ����F�C���2Fh��i���{.�s^�B�'={F	�������lѸ&V����-���^c4�>G���SB�y�5&�$�X`�p�BZ[��5#`$BVS/~��8���g ���FdDR��좃��o�R=���?�a�L�1��4�:q\�bd1� [z��8^ˁO�����n4�Ju>LK�<v