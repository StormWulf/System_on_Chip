XlxV64EB    750e    17c0�l,����o�肓�ǈD���qw�фͪǇ�Nޅ�\�K��k�g���n�ꔣ�H�Ff4}
�P�b;���e���U+�L�8�ϭ�Sj��~��m��^Mo�D|V�COds��1���m/{��cFźR��'|�sLx��ޕ���&}3.r�w���2�s���j�k�`Bˊ��
���!�L�%.c��k4�A�t���Fn;��
���b׽��@��f}�H��ւ��6��O��h�M1��yj��F���Ʃ/l����hڜF���k�h��;�
�eB��)��טU΢�f�����|	�p�@�@�R;Y��a��ߋT�HW�Kl �z�2���o@�,�����rv�b����*8�L�*���~ZB�$�Oj�o�y?0�hR����`� �������p���ؓS��Ê?��LNP,=U��؇%�G�&Q�Mz'��b�3d< ����3)�X������y��|}�(�Έ�}���S�7�����<Y�ɷ&˵C��\�NVX������Θ���~R8
�B�?��2»�cX�5�C_��b��|����p��UCY���n�qؙ�e�&�c�}�=]�t\��{<x��������YA�� �F�9��{V��Te�&j�в�@���*k������,_����ԣ+}�!�'Kvm��7#@ٹ|��+Ü,��V藅t�TE/'�I)�d�:��V��s��v{��u�a��\��GDU�q��bީ�j���w��S�ҒC~�	Z�W�g��0���gp �͖��7�5�ۆ��6��f/��J��?bm(ʈ��ƍ����ǌ�|kˌa�b���]�$j|x׺Pw�|Q>�����y�G$�k�������@j�8���u�����0R�e�)���7�+� 5s���l�#�|5G�Ď9���Q�u�7�Ua�8�C/��g+hy<dA�B�K�1�=�0�/Q3�p;/���x	0S�YQ�qyK�L��ѳ�8&��t&qβ+5�d�\!=��J*8�QjdN^��H/��Њ�U��mm[�T�*�����2ϿDs*{���#�4ۖ(z����'�K���"FL�G'K��L����[��袘o�w�`;��i�}�X�]��l��gu>͜|���H���㾉M��]�|����y����37��l�����������F�$���/�^f-H�������"@_o�>.g��z��-��+��߇Ԩ�K	���M[M��dp ��'�\�]z�b��l�(�̾��%@���)��$K;�X�)�!|��8r$6�@�?Ww��jJR1�_�$�@�1�T	�?+9L�g�+�o�8ZH����s�<���Á�&����D'�CŹ'�����1�Y�y��@qIJB���/�xW�W�|� ���/�)y����K�Xˡ�{�;EghS������`�V�����c�B;�fn)����p�r�Fl�cU�B$Y�z~���2J<3�����}3>c��"�P>��<HW����a}�0!�\-�0ʫ-�t�������g��u��{r�LC����sR3�������z ���!��"5F��S�!�,����K��O�� B��$��3�_�!.}S4�,�L� I%�/�g����㵛�P��3Vf$Vf��E%1:$��Q���`9I��)n���oq��4X����]Γ|�2h��9�]n�d9.u��Z�U��ԓ�nKY�R�KO��ͅK����B�w�}x|��������hd��
� I[J��<���/2��5Z���W�2a!.��)A)�2w�2��ohW�T[�P� S!Az���H.�-T��)LCN�4�w�M?��0�;�%ʇ��֊6�NV�8�k 0< ªzƊTT�IQ��Es����V
;m�Ă����u�3����+���7JΞ+@�9���R�HjP+N����w�NU��iș��O�/�*�	����R�faH�ض���p6�p������I�� D=��%A��4�/�"]� �o����&��<�E� �{8��s�('>�l���ޣ��Z��r��8��������H�i(P������ѐt�R�B��L�Fg�S+?�!Z�	\rLX<�B�����1�OO~���C�/��(�:eE��u(�ী;Y x�-n����qz�h:���f��K��=aJ�M}ם�y��P=�}7'^X�Σ�!��U2��*!�ٞ SBТ�@�gq-BE���J����ɽ���?s�X~G�D�߰�3�P=�&��vB�z�!����A�l�a�}\Y=>{c��1�]�Z��Oª���i�]&��ŗ�
tL�p��ʇ��h����J�:�<= �%BTIگ,�)8EX{|yΪ���=t��u�*����@{snkμ8ì��^~rh�bO��U���AM}h���7��<�|�+�+��s$��`?x�F�;�X���g��̗���#��#цe�_s#9""��.d�[j;��E^t.�1&���Ʌ�FF�D_�C���-��k������O+,��R�1������o#l��q^��VG��H�Aܛ6��+֜����	.#�N��'G(�7�S�I.�@����������6#�3�O��a�	��w-xM0)������Wlܯ��s2Jy�:����,��� ��P���uy�uebqSf�?��[�[d����ӷ�Y<Q����&\.�5`2�{5'T/�5�t�ٛ�f%^��f�K�QAOpu.���t�S)��૏.�X���W�1���㒞I^�0J]��� '��=zݛ�0���>2�Q�wʊ���v�ڧ��#�w���gfv�yBV�z{2��+��OR���=]C�����#�Ǧ��� c1缨��K���E�)���xX
������"H��7��Xc�%�l�BYP��b�Չ�6"O
�g_L�_ ���𛁆A���Q�fp��q#(�X�ܳ�A�񑺌Y}Sk�/��,7leAː�^���$$��g$q��w���Wqx9�Μ�fd�S)߻-W�Y,�����FQ_�a{��ox��;�3��y+ 6d�҈�\��۰��t"��X�%'����Oe`�c�@C�vdRW�)�O+��S&�������!�t^����
���dۍp,LD�Ph�8r��8V�G��e�&��ۼ�?� ȣ3��Q�S��k�+i��C����8�w��7&}��3�ke���⍲�K���9��Y���pS+�ڲO��BN��A|q��;0����4�%��+��Ri�G�����M�l�,���l���l�lM��{v��A+c����K��	�~�o�3�9,�*�-���!�s`nn-ӊ-?���E\ȎHctY�1@�х��r Ϳ���ϙaA-��$��΅|,�,Gz�dQ͞�M޳���<�;+� �� ��A.?$S� �����,���Ǝ�be�x��a�u���D������\��kBE�����C���[w}�GQ�]�p���2��e�<�`� QL�@N�#HX����x��IĹ�U���PԤ�t��#��M%"��
�-��ݧ|H�
�r<�q��/l�C��Y�b�<dl�g�η%��i߼��W�~���Ol:�#3t;޺�/U��O��qV�L.�ԝ=����n��(��+�t<�:�lr���t�1�Z���:WpOT���N�$R�uZ����K�t�y�ZW�y���OuƮ2j2sO����T�t�v����e��	�b_���Z�o����K�YN� ��]a�`��yrFM��l"W����v]��'�neq(?}�G�p�?�=W}�Miቱ���K�E��zG~�7(�uz��!�B7H� ���B;t���Q�f�>�B[�tpӞ4�R�f�_�3J��8�GtJ@��ΊS:��ز��	�es�P�#�W�YlKuy���Y�݄�W?(>��D��xbM�-��25��^������#=��p�X��Ř�[�Q�N�r`Bs����W���C�̜.�+���K=���V�s�ʛ�D�ޞ�x/�/��ؙ�N^�y���ʯ��(�E���mwY�W�$��U��<[!+_�.,WW��j�?��\��]A墷G��Dg�.gܱ�05xi	h$���O6m������vJd��A�(r��y����fHM������m��G[�z*b�n������(��  ��Aشx�^(w�~��u2�v�j9v�������ȠiC���K܅�xE�ŵ�/|Jw������u���aQR��Y�C�$Y�T�`��z��Pk�g�,$^NLB�7�	 �q�p����Ć����J9ǱB>TfܰwÇh��4��8-j��"������x@�+0� [j�}�G&=�n��^�]���}G��O3��=zW��#Y��u����� ��?|�H�p-��^�|K0k�vA�Ҧ�-x��9x<����<@]�3�Oh����]"r@��;�p�r�WY�ް.�/�o<���I���:��PY׉���w��XL�"�=T�a�x�+��ǡ�Hd��lK�4�˂?���{wKv��Ե@ق4Bj\_�|D��u�
$�h8%�mPV����V���j�do\ڀ���:��_��qj����Z���:�\���R�4��-�1ȸdN�v�,?r��5��[��;氲��K�{y�^JID0i���>�u#�F��g@��ӂDgu�+�~��x�&2���J�{�'GRn���"=��~������o;��̭�����#��Dk��q��'`��e�ǤRH){�u��9
����n���q�,�kI�'H-7���J%�z�зR���乷�������Q}��*�}����d^!��l�GJ�r�T妒�v��.�4��4.�Q<g�L��	�i����q���?u�G��o��UD1�e: <�/WF���7V��s?�b$ہ֗��i��咇�	2N���n����؈�ĻA*��ѭ	�&!N2Ge�&Sd�p(|�x�G�Jq�آ��/+���\p\(9���]����Ѕ�?>2�)���H��q���n�{���l:̠J>��L�C����h
�8��� ��B��w���Ca�,�;}��ܪ��)@�*N�~0`WƦi(���Ѫ@D��7���m�z@�ո�o�� R͛j�u{|���3�P�)�4��%D\rE_��=�����y㙳�CI�MK�?�,\*b.��g�V�_��s��cٯ�������^�PU�'Ŭ-1�gU���3,\$��A�x���W�WP\����}P����??�༕���4�(2~�|�R-&���~!W�\Mj���O���w�C����R�i�P9@ �ɽ�rD7�ܫl-�;Z�ڔ^n��<p#P�q`���F���(��K��f��ٓ���8	|~a�����'��e3�a�$$\P��5}��q�2��>v9_��bB�˱�A�`�۳n%��:�&��O�O<a��`�6R��V�:�o/ϽW�,�M!�ǛM$��l^'m!{*ॱ~�����{M�8p�17�A?��WJ��ĕ0<q�.y_}2)�h��"���(��!m��}��½�`�
�dku�4󝝉�q@�~Ȫ���ؽƇ�C��J*Ũ��_^B��(�|Ծ\L�Ntp9�W�M��&jt�lx���e �q��M?:(��>�NP�\��|Bi�K	h+0���O�H�Q#�h���!�c�X!��?'��]��8[�a���a�#~5�j	b#'#e�ȅ�k��m����(WM��3
�v���ɹч�p�׿�yH���vDw�c�g�=*�� Ό�R_���1gP����~�&cL
����U�+ȰG�`��W,kC�4�ɱ_�Kf<l�_ڂ�"q*MoaM�����CO��{�V�x���zZ�"�+�\�\�1c��CʣB/����n���F�a�fo\ㆩ��%SAI>�a1�