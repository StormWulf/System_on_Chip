XlxV64EB    56d8    13d0�Q�Xn���ǠjL�u�T-i.H�0;�a�'�f��ћ�Dm�t���#��Pq7��	���ž� !���x��;4P�Q�c�5pQ#+�6�t�Ї c�F�;y{u�i�&`� �I������e���	:,e�Qn�M��(�"����|p�{�-���>�쀽�Q$t��a���q�-~RP����N2���!�%��1�I���Y�9������:=ԧv|q����I� ���K<5U.1� )����K#h�
�hYk�όR~�x�J��`F��2��w����Q��� Z}Y�|����O�W��Q��=^ ���b�L�f�놠�?�?�_���"�U��B�e}n�~@`����12���"/�)ݨ�"�'oeWB�pw
vhid �N6ن�'�W`�Ù96���U�>c����ռ^�L������N򴽄ػH���*�A*E��=PL�N�;[EQNP��$i�"��َs]�1��"�m��6&�a�(usl_f���GK�o����9W�������cc���`�5����1�]�z�S�	ɩ�=$]d��p�x�9�t#������ǳ:�\��8exK�ۼ(N���W�gK�;,���-�Ë�_!�!�J��0��s�X��,�C�c�Q�I�Q��#tr�D6s�_Jw�Tw�ϔ^�#�<��N:A8z���0stD ��U�;bt�`�t�EF�����/�ȿƧ�L/B1]0��8:��(�: ��x��V�V��� ��5�ɱfK��N�����`[��b<D���ɫ��j�c�ٟ�1ɘQc��(��q�S���N?���q�	m���e7�hIl�.��SWא�\GtOd�g�d���°)�W���"�[�C\A���AY�����*=�V��Е�B�	a:��z�-�8����9�BN�̑�o@7V�!{�ơ����D�I�Ib�L/����	��z��ŏҸ�e���x�]�&@��ᅨ�kL���}��:=o�H�F��'|d�C��I:�b{���q*�R��������@��^׬(���}Gy-����99:���n�lD4`ō�l��f�C�r��GǗ�[}�!	\\7�����؋�Q؄/v�� x`�0��
�z{��E�be���B�M'���4�* ��^r[��� �!�bB�Ǿ�M����F�]�����#�YzL������Z�.��%��}�#%�㕜�f7G��͝�j$�h��t�5�9�K��v�{-�8�
M��>C���Hz^��um2���g�2z:��xk�������C*?)瞏��)�Z���ny�����ym��T�~Y�=��u���X���	����(���<-َR7��y[E��_Q�p����q�t_%�<{��O->?��r9х�$��ʁ���;���.���%��מ����Ac��l��&�b&�<������O�&$"p	Yz፯�C���{��������ڻD���[�0<Z�>BBبܞv�c���~�J�jN�u:#��	a_&�|q�Ĭ�5�+��wHy�_T�#�c0�K����� ��{��&���[]�_?!W�U��(P�j4�8��'���5���r�14=�>}]�c
��n���P7p�)h]G;9�S�� E���KioM�-*�c���������k�JYC����񒏋A��~�uf��P���h��ހ:,�*డI3��C�46�]���
|��0��,���ܠ�.�7�6�����u������2S��ere�F��J�D.��hj��S5+���,q�q"-�R�z�J��A>ʭTжI��"E��1�����l�_��� rdD�\oޝ$����~H�0�<|�θ������	SD���>/X�=a~�� {�ĭ���N:*"W}n�F MθF��8���5�XUF�C�"i#��ү4BF��c��~ڈ�;�L3����~\�%��qqTLعF��֣���-U��/��3��W�ҙ���>᝷4�v����P�R	��`��QvX\��*X��s�͆y����w��v�k+k@�9% yG�φ:ɽ��4~#�!���	�\���ې�:@΅���W�u:)�/� :���/������Id���(�/h8�}�"`���J�	%̗�����49�B��� FC��7w�]��<9�2��P�Ѥ�)&�\\�7����n�n�:�`2d]��J��:�bV5b���W]pރS���(Ԡ��� U�RL�>V_�F�a�!�����0�E��i�i�-�!��g��q֞�AS�������0�������#�;9�ַA�i]�������Q��)�"Ef��P��ڹG|��ZϴɃ=�B���Ʊ
��*�܊�l���{'�-�[܄(ȟ:=E�_Y`Sh�L1����&��n�G��6�~9ڼkȾ *����*x�h�s��wWٶ�%<�!���L���3C���Dy@������s,M���6���׻�^V$�[T��%���E`$�ŭ���r��֯�T-F s�L�8JN�Y��P�<�8�]�7�a������F�zb��������!��$���'g�!4>O�]f�2I�^:Q��o��M:JN���Itg���7��2�0�m�R�I�sV����.W�dp��0�²Y��Hr\�I�f?�3��G$I�� sC䁘_n�ܴ?��A���(��b�����J}/N�.^v�'�C	%wY�~�F�?�,ޓNjH2�lM������	 ��J~,�Y3j ��0��g���u"Wj��0񢎲T"���>^.�Ag0��j�G���	v�ݚ�����t+�I�`c�O@����R~s���jW��ʧSE�����~A�Do|Iu��y�䛔�s_��3��-@A��=|+J�jމ厀����R�e�_�R#{��Ŝ#���
�{~�9���3����v��*q+���G�"
�/��~B��d�'HorR�;�j��$�=����
�0wtwXP*�$�m�1@j{�0r�e@if��󳾧kݫc�p�:����a�)u��fc�넜�3�k�2��"��~rl���b�X�->P��j�<	�о͚��~�a��N���{8��솓��� �G�b�I�I���<�[�����Ѕz`I6�U:ֽ��+}J��0�J]��ƈP2KƝ�f���3��^>����J%S�r�?�s��}�1G�,��ٛ?;�b��:߈5�r���	�ׂf8�� �?#Y]�5!WP���{�-s��Uo�PC)�{�y��ږ���
H����
���\���(�����{��eS��Q�.������k,���&���"1B�g[��%���c|������n+k���z�x��M�����Z������7vuhe1#Rhc;d�[�x�.��s���?�L�s�}��m����s�N0C~6��U:�a�V�w�l�b3P!D��fy�>z��;#[��]�1��b�s-LH(�H�����C�$�J�k�Mݛm��!(�R� .i�E�2�L\%���9�����2均�s�\2�W�u3yJ�����X�2ط�8V?�ѻ��^+U��v'a|�b��M��$=�����A+�2׹X6��&C���%T�(�q5j�ƶv7	nÐQ��7��_�В��/O ]w�X��$,@�+�`8�&�(Y�s��ZrA��y����?�R��ǟ�aXaB� �U���u��5��)�Yr��);�y��R�6��W�5��������/#,�� ���O5�����\����&Z+I"y��&tf�m�PG��W۟|l��D���L��BFW��1�?vMoS�l�BX�~��r�T�@}�'ǹ�g{;�邔K�>Ω�af�a����; � �jhh��zD����޳ � �j"��R�ܾ�N�e��Xy� <��jC���F;B��1-;䗴�X��M���NcXJ#J�|q (2��Ţd��#�<X,������H�>���+��]���<}��3R~��tfZ�Mھ�r{�A����LI�癥{5��A��j�q�����@L/�Ӊ%��9j��b*,/��|n��aZ�ّy�A���[1��oޯ�a�K����KN'�s*#��n�@Aw��kn__���f!����l؜gA�=�F}
�,�jjk�I2�
��C�2��jZm�MVB�z���r��G�O�⸖�y'��(ާ�ث�о󢻄j=D�lE+�h��u�%�l�� ElOP:���ɶ��S_ΕK��mm)�� �u���L�rf�2g3H��E[�5�BfCtn�b;�A5:���aT�&�1�W-T�0ZR*BU2o�u��a%7-��t�ޣ�>Կ�����3�LT':J3Ҵ����i*1�p�N��hC�!�'��|�&}�WD������uע%����%�,52g�6r��9��/��I���v�9h r�S����%侲�F�.�6����)4H�lQ�o��h�Y="�^��$I���!Iم{L���̗�P����w캩��.��v�U���� ��R��Rq*@�#|*o�\FO�jr|y��#]о�2]�bCv�ݤ�[����l�8�]�C`�Б��òe��i~P��x�ً�1LOp�V`�k~�'k�xu+[m2��	&���� 
Z@-�؆�D�N��4�")�����iT{$�:��5$�%f'E߰����P�8�̰S��ƎAB{���&�8��E�\�7���*��b�.��H D\�C�=�u��s �eQ@���R�������B!^��3&K��O���;NCR�Ex� i�(�'�����GB�����S�oҐ쏰��L��t��u}v�{��|�&�m���߾SŽ�\P��Fmzw#z'���E�][��M(qo���e&��>RG�.�^�c~�z�j���S�{����rMm�\Ɵ���~쓫 �q��#.&��P!}�{�`]�HVq|��d��T�]�9�sNHs�S