XlxV64EB    2a70     cf0<`�0[�����i�=?`GWKk���uQj��Z�e9��r0�%o�y��h�S�|MN����`?��($�%t�fؑ�D���{�U�e'aSx��,��*R�O��@��*�~[�/��sY�=ص���V%�.�GI���� 0���\�߷����ۃ2\<S����a���y|4�B<fg���T���x&�b�#?�7*a�rB$��j�n��t�?�m���gO�6�V^ؚ(u��n�g�"z�G��)�� �����g������܋���g�6dߩ8+��I�q�u����^!y����9�;�(��̌�<��M^ꨟY�8^�#�J�;v��f����ΟH�`�:���P���E�y\��f9�#j,gT�@B�թ'�m��[.��U�Tf�U1�aA���"��P&�Nz=%q2"��{��ne�K�b's�5Ғ2!ɅCq��K�o{�"z�^k��MgL~IK�'��`�P�۩�*y�Kmx�-B�R�b	Fa(��]�ɝ�ZÛg������h��?��,3�Oؓ�a�Ť��|1��߿��z��t��y��7ZB/��̹�Ztu!��������l�	�v"4<sX!�c�fxV�,ڨN�\>1�����-f)�Vg{�^k L��kd��)��ѣ��g����kV!�Hv_Pu?՚��S�$d4pNh/�f!%����I��WxotK�,���<��	��A�4
����h�yb}�����aX��ٽ���7�c����Swu��p���\@P�I�G"J�6p�`��{����p���:�]�Bh�i��7.+�b0����H	ݭ-)s(
͑��2)n�?Ͷ�`1�$eR�����I�MU#�i����|q�GK-�>��
J�6]D5y���:�Ei?�n���9�V�J8>�~X��g~����Iw�cc2%�~u�~�n� �w��z��JP�S�M�-ා
�w1\ϴ�)]o�oNLd5�2��~��0��ɊQ��WK�M�0�?{�����OzDc`�=n�f8��C���.w� �Y�!d*��/��f?)Q�bT7����$x��s�A��]�Ӱ5����a���$��{,��ͅ!Y�g�v�&����`LP(O�}��_���D�h_``y�Yu��c�s&�>�ƽ�8�4P�3��=6V<�u݄���0I�w=�E��B�$�v.�n�@��KT7��A�Ь��yz"�T����&
 N�t�b�p��}�=ts{�˅;�T�ɕ{����/Qq�2�?�v�4��U~
�r�mKy����1bj��k�m��,cdz�o��<n��0�U���qrY�O��r�Z�{=��~���pW�zXO0�A~-��{=K�tZ�x)M�b��4����X�؄2�$�+$����@>�F��}8��`�'k���F�Ff��8����gv�/],A�-qK��{�������@������}�^��6�p���WǷ:�7 �WǺc����ϕW�
,i�QD�]��p�����Σ+Gm-QC�'�NI���	�*���.�8o�� �E=���z��SG�<�+�n�n�7e�%��� r鍮x�&�؉R��OaT�`�vQ�bv�!��N��=����D���f'J��4� ��@Hؾ��o���NC�(������V�#�r�`����sը����pu�[��o&����>p�n��А6I农�� |��+Ku���w�ؖ�2ٽU
��u�E�9x-'�h�[��G��1f��˲�R���+��
���O1h��^ ��Ŕ��A"�ַu�[��(4��yx��;Y03���1fL!TO>�Ks4����=o��mP�Z�T��%�(������i��ĲM���z�ϭ>E�*�m\	�w� HE���!8�/��*��L�����a�[���8'�Bd�!BG�b���]���dy�P�q\�\�8�����#6 oc�����ы�cp�A�c`�x��8������\�0�����(Q>
���c�Q����5�{p��<+�A���K�v�[��Nt x�,'���ߠ|�.�x��w�	1�*�5���[�~��D�+��pB����]�Yɰ�Kti*�^	�1a �n����ުMrL,��a0�鐛|(����G	�*�\�������,mӘ�Y�����אָ�*JX� �Z�}U(3��5�bA��y49���Ki�ؼ�-ɶ���C�'	��ۋ�)ᘳJ�x"�L����Fe\�?!5�����~:����T��6i��N��i��ì׺{�U-*�Gg�̐�oL'߄*�=�I�ND*�t�� h���s�f:)г�ڮ��}E�(J����M�-4��]è��¦�o]�v�	�ٰu������,����-��vw�gS�fAMu��[�i��4f�wjA� �ݑ|P��>Z�͆S�7/.�ӜT`i8閼:����������o�v7�u����!����T'����(�b�ƣ$u����^�SYV���p�W���j�1���vL�S�ۗ�F"�\�/ wd�h޸�p��<1+�A�X�Lɾ���i��/�6{��e>>��hT@NMR�U
s/A���D�62,��!��g��>� ��������8��6�;J�y2��gˮ�f�y*
�5
f}�3һ�r���vF��&x�JG&3SDQk+`�(y�|��Ā&g�*2W$2e�#����i��fl��~�x�*��|��0v���N �ꙭρ�$�1F�E�n{g�;w#�[\�H���7�Q�P��jq�E"��ٿVّ�u��������d)� ^���>�^!�G(5frf��|�𧃼e��ac��,�0Y#����7�S�|j}�R�OAǩ^>�깰��Q�Q�L�u�6ـʱ���̾Mr�}D���hf�R��U�e4uSp�V&����@�����Q�N���ePZ�����G�+2��1��b8/̹Y6��ۘ�"�{{�i�:4�ϱk_ﵫ��m��C*=4�,�`��^�h��)�@y��f���W��N��ѳ��g��b��v6�]�����i,q
v�5��O���x�ť֎����_,�!=����*�~�5l����h�09}��쑤\/�E�|��zQ6x�\!�G_c���U�7�k� ��o��1gT��-�nxx+�.h �J˵�?���l����{!���C����%��zŜ��5t5qZu��'<���W�I�jA�w#�e	X�&��/���ШBv����H��e~_�]vk����f�d���h���%��CM�*�5g
/u��хP��