XlxV64EB    b70e    1bd0p��B���@Wa�L��y�	��V�ӓE��d�x�s�iV��XR�	]�O���`��ˤkY���"LJ���xC��FL�5{��9<�B~'�\,y77��8�	1���1nAO0藗�<I`���&ߔcr"�*8!㉖��b~RdgO}���v��F���FWXڙ���*�G�-��e�F�<�˥�<>���n��;���|2����i�m�\��	�����X����������I�s���*OCp����n4��\�F��`XG�H.�$f/��c���aU�	%�P�Y���g��q#��a���ƗֻX�qY��7ea ��������G^��C��2�m��7�A���y6m�^�۞`5������k���Ѥ##���P���נ�ņ)E��������ӻ�){p�gDNe#&9j���PQ~gL0��t��+�,"����O�"r�(gG��5qև���'�N����dB�:�$�XkgO�M�&s��/����(��P�æ��{�#��GN{�/��Y�Nn>}�����l�p�!I�H8��̈́�_���@���PCn��$�2�"�� g&�-���g�:O|������饧�y#f����&R᳞�5JC9#!m��PE)&z�E�$z�'���H��$sr-x���zx5��f�'���#(h���e�@�	J(�jG۝q�ك�y��.Ƨ�>�̭��w*�|�+6�wG*��C��M�6u�~���!�
ռxM�����*.��a�U��b#��/��W�5y…���Y��$F6��-&�������|�|�l.����;H
�������0ŉ� ~�賛��*����<���'�f1V���rMo��N��H��4r�X�&�z�m)�`�#7T�c�i�wVPp�o_�l����M��h�t~�x�شk�Nو��^}l�+?6�&r	Ex�b4v����a���PG��e�mv�}���z����� ĦX��L�zIF�~�z�G�}M�qQgD�E�-��YN�	s1͢qE��C`*���k�-��y ��qi��!��O��IV�5�_=�I�y�Zc F�䩪�X��$��TӲ��2�}	�{z���c�2E{��O�,��ׂ�	�Xp��ˋ�GH
�3{C�a&��;e�C�n�+6	hG��.���~�\��!��]a�~I�'��|_ �H����ȡ�X���ϗ\�su��6�3(��Sb&NF.ߧ'��VS۪&��J:D�^�'X=2k��9�1D"�=�~Q&�Xa��BE2��)��x9^���=�jS	�D}�hX=�ʉ�$~����J'����7������5)�m���n�W_�m��XX��1b@_Kq̰�"�E��[g�U'Z�첗��z��Ш��!}���]�T3܁T>���`t�P�'x��Yg�����acR7����::<�{i�Sb����|O�����:��|��B��?��u߆i���a����|l�jb�&�z�+ۖw��I|ݒ�K$�j٘ז
Ѯ���jbaQ��9��A�����כ��E�t�<i�g���S���V2��h{)�H�$9��q�<�e!����*#+���c�� �62����s�=�3[�9�Rua�4~.�X�;I5�{�!J�SDboc�x6�H��׌�=���#VD���>'k������x-��0鴖�w6ό��'ޞ��#�������.�%ՠj,M>*�!DDl`d��g����<�L�'h�,�[����(b�Y?����B���b �{[1�n2̞��m(ߨN���晰��Y��I
�.��QMp�V.���h���r(���������뎕�����=��3y�F!d��4�'՛U��O�2�~�W�@d ����=g}:���t�X)��ػ�~VC�Wڽ�� c��/�G%�&�4�J�bu�K����(/���t(s��oJSM�F�z�_,ņgs�E_�`O����S�Ǎ%Tft)�w^�?"`Sȫ�U�:v��#k��6�O�M��k:����k�b��졦N��9���l[z(�O��=�.Hq�)�z��/�/#�t��l��Hbm�mMؿ�Ǹ�H�j��ʎ�d��i$�R��j��õ@d�1�mZc�x| ���B�+T���
L��q��ǚ6��5UG����&��/�I��5u��:+��*к���Cb��<��sK�8�E��"�!&4n���No����C[�0�Y�	�l�i*�Y�����z��>oPv���I��,>=�r��[��o��p��+b�>~�WLp<C�IQ�dڪ���x�q�?W�U��]+sz�SA���7/ 2,��i)K�`s1D(�p*F� eX����&M)5&�.�,�s�q��o^�%v"hm��`�`gM?�%�����J�)���/f���������e'����6�2Q7�'s�mm-��)�����=|�k�r���	�&��[ksC����B�/���S�G���F�G�;���e_"7mB��H���{�q	������y��T�H�Ҿ@�\24ew�U�~|sW�^�N?�����o�T�)��ɲ���Ko��#g�+�5�!�e�k�_�o!���盕�a�nd�?�d�"U? �e�f���.���t�*���c0C��VT�Ü�l��&9���U;�5�����sJ��vg�̻����)0>�f�oLh���+Q|/�m=�1����ZY��k��8����+�����&k�ŦwMKQk�xU��ρS��Ph>��uX �zm1�L_`L��6Z-�Q��1��O�b7h��������F�	}e�s͑���A�yaO��K�wi��<q��i�:ߋ.g��&���[�I�6�)zu��yO@�w�F����m�y�,��%1�^*����Y�uq.�*� �A��1I�O�MQ��P�?~����#���OqM��M�u�n�8Ё�����j��D�t�Ļ�${��ߎi����H2epら�sT�`7�k�I;�,�g_��AwK�EF�L(����	(��_#*�艨�ww��M��3��G���<Ze1�k�__�}$@�B^����o���$Q����x�˝�x���4��wʖ�r�����p��<�Duu@SHl�&,s�>m��Y#� ԃ��xڥ��LGn'UIVy� �����
h;��9��U��#Ќ�mS!HM|Gk�{t#}d�e�����$��I�2��V8N�Tr��v_���K��y��q��4OaC��N�
m �+�g�s�YS{�,�����|g��ߟ��&U�uy��p��;-�Xg�j�/�N_+-��gP1w��.&��,�#��v���B����! �e��	�5�?��K`�I��~�T�6=u���]y��va�Zu�G�

�saH��O���"-.�"�Ս��j�e?���-����q\�&���� i�[f���s�3_G��P�ӣq4�y:�\�^�^��#n�c�f�<;�#E�RQ�����+<��}�@���]"���!h`� ;�1������!�;;�$��R�א&/j�ن��>������ H�P������U�D.L�QrN��ا��牸qr�
&�-U�����j�]�M�Y�|uM <�Zkߞ�3x�θ�V췃P7�һק/z�)"�V]ӂ��ې8LK��V�)����������+� d�~��������.���v�s�pc�3H!h�5�t��[n="��KZ���RxR��8e^E#V�E`�����QS$L���2.t�����rs}N�0,�G�9� ZN���L����@~���ϲ�U�*�g����%�G��Vv��f�v�X�N�#LL����0�̔�?C2J��jw�f�Zbf�a+���]�.����Ǯ4�����i�0�N� ���e�`Ԯ�"A<N&�ӁE$�Ø&�Ks��O�E���DH@�3K=wt�3��\+�١�.���I�%	e���09�Dn�=\�u �
ǦĀ��]mzr������o%,�.��ӿ�-�z��[%R��+Ék��,(p2/)]�����G���%��g�۴�Սo� �UH=�ϋZ�T��'�$�9�6��}�(�4ѡ�*+������5ޒ��	��Ω}a*u�g�%w
c{��"��?Gz�=����w��X�y^Q���Jֈ]�7E����M`On�s-�T v�
��#(^kw��K'�����|�.��(��r�H�2�GDXZZ��^ �Ɋ�ߵ�=3G�SK� Y���2��`����?N�~7G9�c��(d���Aؒ?�*	9����mn=�fK<�Y~[oDNy�2��9"P�w�@�`���a������oq_���w��i�E�}��5��D�uQ����.�����O�5�L%(�N%�S������D͐۬�j�R�7ܜ��df��H8}(ѥ�����Y�F+����ꪎ�q\Y�U�MLR�Ln[sb��g*���Ѻ@������;��qy�d)����=��e��lt؎`�D��(��d�k�E�d�:��(�!V�V�R�E6�����\�1���Q7bS��oA���MR���9���#����U�n��zҩ���J��=k��������`�y'X�8�����p� d]����/�P':E���Dw�A�3$��)Γ����*����ƕ+�����t�l�(�V'�1/�X�gm{�'J� �C6o�o����w���^Ⱁխ+�"�G3$�6�W�Z�-D�<K�ʒ:}��ܬ��y�oqY�'����a�QpL��ߒ����M��@]�X?�?L_�>ش\�g�(S�KT.Ä�R��Č��S�X�B�|^�?��ԯ=
����)/^؄g>�i��������4�^s "��0V>���5����OO�b����G�dncL�ݶ1܃�C8��w�`|#��H�?\�%D���܉$�?�V�(�p?�j��}l�|Y�pS��)��4��e��w�9�'}�S^��c���k)�!��MS�Cu����!pS#-&��ۈ�7��
q �p��0��YuIE)�+<;���AC	`a�
"@DĂ���Ő��Tt��u�3�VKoڲ�(d�Ǽ�Gp��{!BI���L�(��������&ʷ)Ė4�>��҇����|� Ű��/����g��:5�e�e��U��O�[ފ�ݦ�y_Kv��DIмĉ"���P��W5����&�s+R���H��be��fd�wH�������#��s�2m豟��hݲC�4S�^�:6DY�Lq���pU��š�XY��S�f|��հCK�P���ա��o���GбK�a�4��@��8E���/"����P#N��9�M9�(Ɂ(D>��$4+o0 K�>�s] �T�)�B�8mm������$�V풩��{"G9�8A�� "���.�����cm���VEf�q�y�i�Hӣ�J���PHt�S��27�B��O� ��w�r�i	��Z�xX�5��7X����YU]���uo̴�X����l\n�䏪�L��U�(�w� � N��Ir�:�ȊBw ڛ���1������Mz����m��Ny5� LYM���#�;=r=+��|����^I��=�ޭ�h�/$]�Y��JMX��:k�f���Q,r���+FGE�����7��l�qU�e�n�̋�K��rQ����f�����C!��ܕoO%��O���%َ	#6�����.9�]E����� ��֔���'�LT��_���V2��ߚ6m�*\a%��p#w�%<h���k�6&#�(�+Х����뙤9�Г)�`�*�t��m�q<�4�ئ��F�����n\O��:�s�_&��&�i���_��7O�����6IsR�>γ�Y�}�d|����zHV��d�qOA	�� ��.(72�����g�&�H�|�ٰ\,K�0�{Ӏ�{Ùǿ���)^�0nKԣ��ز�2�}�֪�g;I�G{E�ݢ��zO����C��'�]_�J�M���4is�qonK,��-�'���\H��l�^W���L�{"/	�U��gj1�7��H/��gI���Ƹ�V��M}��D�t�"H/&Fs<9�c��b������Mh7�V[ ��#�#j�~)�ɳ�����Pʡ%&�ŝ��su`��G�H~9M:�ꔮ"�3uJC��#��Y �.fV�&�h>��� � ѼKH�[�YI�aW5�D���{�T�Cog�P���>o9T�g�fk+���:neGEV֎m9>$%Vh>Pyٰ߬bu��i{ �ܵ�_�U��CS>VWh���%>�rIrOU#N�9r�Iz��Nma=� �a
©�Zg��=�� M���C�1#�T $�d�V��������.M�#"�StS�e���w�Hw����(=����=Z���{S��ȎT_]@���ؖI�*�q�����S~�H�^�AS?-���}�*H�P(/�w��A�< ��m���.��X���s-P;��A��O�D����,Q]�&1/��[n���N�>_��f����h�h��Q���!�s�	�*̽�f�����W�t��H{�Ej�n�$�M�*vgh�.��ֲ�E�R�񷠈45�^j���<��g
w�x,�$��Yq�����<�����������ڳg��¾��9'5	����V��i�ĒL�l���QI%zX�'�Mp��	/'�؞йڽ�"E�$!*ȸ�m^[S�O��I4�P됷�[��Y~�8fؿR���.z΃��><@�T��H{��OZ���i�N����P���t�K�ޘVy�T"&L�/����D��3Tͧʗ�面�LpI�!��XF�٢��x�i���6�|��8!Ϝ�f���*(.�E�z�t�//�q�>��,�� ���Gf�É��9Z�-A^���^�27=;��y�B=7f��}ܬ��f���~���]�biҀ=b�ӗ�K�Z�ᆌ�p�&^V�d�ʝl#X�)�`�RN1�t[5�{믷�Q(r[��aR�ϴc�aԱY��p\)�1\̎\a(�x�.3��'�Z�9�i�)q�A鿄E