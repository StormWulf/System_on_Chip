XlxV64EB    1d20     9f0#I�a6|OX�w-���r�M'�f��ЭfpG�} �����Mj>�A��pgA���&��(���Wss�wCS �x�|kb��U;�.~�]-JF4=_o:XD��7�,�+�,b  ��I�}Fѐ%��i9.q����N�!?��.�Gb�8Q�\��3��)Y}B�[��8SA�A�"��5=h~���.�zS�]�2��x�\�l 	;v�D�.��'za��e��0 k���Qϳ�����M{	��v����pb�jE8.A1$~)�����$�
?^��8�3�:CP��L�1K&��5W̹�8Dԫx��P���]cC�{���|@q (C=?��IH�]t�}f~"��&���'>O*����UEZ�~�r��)�Epr?W�uV�x����,��ޟ/&S���}��DX�Y��o�k�p�W�	�n�jh+�;�����3;�L6�q�Y�b�/�s���RX�f��w��aMie4\�/xiH����0w��Y�x�$g0_�?�Z/�;��H)�-1�O�����<�Y�"�0�,���'�WN�M����ti���L���ޙ��t�v�O���@DֺqI}s�L-����?)�טs�"��LA������#���skE��d�q����'%��������@ Jm|��f�Wҹ�o/"тNk�64�.������l��K��W�4�ub��Ś��\���v�V;�޷��vnaF��y��/��<�3���AN�M����]5�eK�,YHC#j�d��2��̹ U�����<�i��֍J䱿�ʩET� #=c�d��������Yu�����������T���Ɠ�����H�r �$����H,�O�.N���<xa4g�[������9���]�����kIp�[�y"v�p�-7beͯ�m�%
ˠ�:�706���[�,y��ZR����P5�&�o��k���҆N=)HF����@����mMѧυJ}���%N�B�І�d:b���w qa�v���'��!�u4=ʘ��H��~J}yK��JE^z������ü���x
M\~(����ݷȸ�<�b�A6l$��^bެ}<W�:^�#�S��I&M~p�Ⱦ�k0+O��X��nu�
 ����ը<S~I��_H�3��*ۡ)����h�+Әʦ�ƭ{$�s͵O��«b�\�c5�(�_�����ī	`Ft^�*'�؉��⛴�W��U~�	�t?��	��y,׊
�q63��rΑ�O���D�~	���Ui�$�$͇�e����W�$�8�I�W�l�Ջ�~�Γ�wp��v7�yI��p�� Bx�I7X6@0i�Q6,"�8.�l�鮑3���\H�%-��s��	9@l�Ӫ��*���%�������f|�Ik�=#�&R*42����n{�a�!��T��L���Ad�n����WI��(S$-����&Z�$��1�~nT�L߂���I˃�R��,g��~���w�!g�a�5�i���RNrMpZ"/F5=J�l�CsJO$�r���4b�������u�F��h֧���A�0�qi�l�;�|J�����Z��-�5?���\/*.DA�ؖV�Y)�>��3֢�ha��$K�2�����(b�uL�X�YbZ��]�����M=��O�B��0�c�^�>[lI듎�xsZS�ɳt�T ���6�T�uU�u�ֱ�t_Y�0�@���+I=�*2u��g4�S5�8N��.4] I${ L`
/d�7�a7;ބ3?��Mp���R�H�P\�P�=�Nk�B��:�s]�ѽ�6v��y(˴CV��xm�2̣�b�G$2n��S��b0O��z �0��q��]��a2���hP���yH���c}�q�a���S�(iz)9۹I[��W�;�x��Gl:�����n�i������4�p���N�)�`2�:��t�V0Z�CҲ�l�N4�w��1*z��C��W����Fu4�[|v�i7$��CyI�E�t���v��f@"71�x\C����O`~"���E�����I�m�W!6А�'����&��V����g{:��^s���:�<į�^�u0}��υ�{!I�����>�+�E�.�</֢x���2Cy��8�qe���\�E�����K�ة-�@Z�f�8tr�jUm��^��5P�=�Z���# �v8�7o������Ӌ�y�QI�B|�7�(�� ]��-���_�J�� �/�(x�F��~�*ٱ��g�x�M2g9��ub�ξ�����c�w��Ⱦ`��`ht)ښrL�*�mVӳ��6ՄB��^�7�k���Ks�w�ϯEh�~~���9�B��}rVN��~<�X&B��B{�	Riw�!�=`^Ļ��p0iX�_.������,�j�C[ qG/"p�hi�r��0HG��5�^�c��+�*�K�s��*��X��&[����i���Y������W��ah��W��@���Q��}���q\���U�=rM���if���֬,{4ĢLj6D��������p,���