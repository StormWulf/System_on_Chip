XlxV64EB    15ba     850.�Hf�g�?p:�TB��Er�W�S�;��ti1���+������e#J�̑hw8��R���l�W�27K���P�<��D�LCͅ���m�ӿvdJ��Sg�p�݁�Bꅿl��?}�)���B�K$<��;�z�����~� M|1?��?�d��B�%A˦؜�a0Q؏A"�EޮF� �����l<A^�D�]��C�|zT:��������WTƪ��m��᪺+�;��+��%��1*�P*���u��NN����9�� �D�s%v��B��V�R@V�Z��E�C0|�V0f\��X\7a\Fa��������`�2����ִ^`�&���1���͊�B��Zu��&K�-܋�r�%V�>�i��vO��ә_l�Q�4ȐwOx`��|l��30b�����5�~�y���ʱe�2�-���?wv����"�uVK�}��}z��O��+�`�Oz����R3 �	(���.9�����:h<Q��� `��À]�~+��RǫPYq��|g����悅+�u�n��X�;T5��KQB���_���5�9��ό��C�ҥ;d:uR���m����Ʉtek� ��֠|@�B�rr���l͚�E���@��`:��=�'n_׃�Y�S�����`��
#s`�g��3I&� ��\���d���7���G!������V�9D�{C�.�0��!J���e��J~�W�{��I�_�����/�� ���,�
b�yiط|_��:���(8♇�Բ��s�H�L�F���9�������IF]�/��s;$����hrG7�߽!:)��g荏� {��yc�1�:�ZT��?�{�R):�$x	ۅr��iIS�Y�z4N�^��� n�C��>���Q2�聝�8�r<�G3]�ަ`��x+}v����a<a�����J���YE����'N ��ۚ����'��G|N�m�V�˫�2��p� ����2��L�-��,�W��u��a�����14U�3�厀5mb��Q����f}�eWi�n�{r #a7�����{�]�u?=� �@(�>�g5Z���������c�r���|�T��+��r��]0V��3��fe�I���>��"6{座}�g�oR��e���R���5=E7yϙ$�Dg���b~�|s��/H�	��%h;J��:�8Z�t���S	�����ݛ���yY�S��N���]C�v���`����QZO��fd�M��Gz,�4��K��.O�ÝP�f�-��<���� �F���P��]�-BS���f���g�ךs�s�7]�r8�C��x��E����)C�FL)
��A����_K�7��Al���$w���?�
S�ѱ�+=�=��f8���,i�b�2�]k��eL�����`__w�M�È���s<�x������,�YM�0��Vp*�4�E�j�%���YN�I�&��gb��?�uD6��}pt�Ǜ�@����R1��J�Q�y���T�ԑ\^Pi�O!�?�՝�͎�3�qzM � n�$��9���#޷beP�����'N����[h���<~���+1Z>�7�����S�㊰�p����p�9�/{�x�э֛��OrL�u>mm�|�vg�A��+`\TD�X�:��췀�A�u�H�+OLv.���qK{��B��Z��^�8��E���R�#����t�g�M6�M%h��z�j�n�����c8)�\�S����+#MB��v�h�?�+��q�]���گ`b�2�g7�Z�����,3M�'��t�Ȧ�i�@?�LPg2T�4�26óp=���F��RU���
�1:�;����VWh��0��O�B�ߟ�� ��s�@�8	���fn�#�S�u�G;�t@�qQt�ҵe�v��09jZ��MV�`���yE��N�����S��1�����y�:�����N�b���dg���+�Bܡ?���!l�����R��ytv��k{x[T e�j+�<�e�:Z�T�&�P1_��D�a�6���Bs`E#��yYՁz��{4A��F*��Ӆ��I�?υ��%l�MaFƒ�G�����/�0C8�[v�����K�7�#��S�