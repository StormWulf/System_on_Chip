XlxV64EB    221a     ae0�+�qɗ�5��}���?�9!�Е��/����Π�z~�������z)��ɿ���q��\^t@���D;��Z�l�JD���7%�.�k��f"�L�����U�)�ܦVIc7gMl���aч��#<�3��ŉĂ ɲ>�OU����xN��x����>$����A��\��G���=��jU�8�^�њ�hrd�C��l�̅��&�q�Oc��YLˍ��X���$�%�6u��;�s�FGt���Vk	�[ki���_�z���a�S��"�@!f�H
I���F�Ն�I{b�*A��9`���A�<�s�ժ&�'��xT����+�&hv�u�bIo���ѧu�/�9����Ҡ�%_�=�vV:q	��EY�����)4�4DQ�� pա'�:���禮�����\]A��yC�b4�E	*�������!֢�F���O%��za���B5��5�*m ���zg_�A-Yeeo��?�ccU�IN]Z̡)�9������a�S��_
�j�yo�mI6���V��@��(��f��e��Ǥ�gT�PDx��@~�;U�	"E�CwW��vѺB����|��ru_�,»`���ABQ��L�:]�x_,�9�|�l��f�L][�R�{K�tϖ�v������m~�������Mp% ��뫂v���ͦB�Z�����Ե�~96.��������F���O��B�oX���}GyN�קo��� ��f���(�C��֋nV���c~S���_���L�<�\�-&���&$��7�h�;0NU�iU`[���ʇ�����6?w�E����g�kXj�X�
��*�/�I��+���/J9Z_b04S�!��	aZqr&3�l�щ��f�_��U)�&�/f5��% ��_�M/b�4߽�O:;��IW�V*�A�Z��(d���;Y�a�S�{+�6������&�3�u=$3��Zq9�/%���w�a����3oG�T���0O"_Վ�y�VF��RjBRמ�ݸ�t��ȍ��W���.�pw��r�Uz�*��2/*�NX�&a Pش|Y)�&w��<�v O�T�U�p���܀���tv�����qpZ��S�Adm�4�-�k�m��
�+:�~�氠����aZ��{�b�t1%͙g/�x�������&���V;���pfR-J��5C/���e�KR�5"�ۯd����6������9�L��@�q���V�	cOg���{� <Y�~�3�ߊ��uV��i�]��F%U�e��-�=�SWo��@\�aO�K�<Z�+�l�fL�Af=��=�SF�Q��~�{�E_���O��<I���O�Q[l�ݰKf���r��/�~��v�E3�T���H� Eh��=rӐ�e���]�_vT�r���������@'n�>��mW��<�H�wth�֖�^K���I�_�i�E1�v6�ҿ%'����\�=����ԛt�#e�:�O0�7��9\��	r�j���Ӽ��9ιcgR����h���ku�֊;Ԩ��7P<or��;� �Ą�D͠2)0���4��*���?�a�}��[��ϛƦ����m��1]�k;��t#_�5���I8溭���-����^��t�>{�Oftt+�s3"��N
ڋ
�.*��v�������X��{�*�D�6���k�����~��'�*8wu�������ɪ�*��%�k^�̿�)�/�k�퍸���Q����H����w�Y�{�t�f|���AЌ�����
N!a�k������o����5�{J���]�1���D)�I�nQs���O���/_r{Л��j��>n��৓�8��o�M�S�U��w�3`( fN�}�H���R$�]�2�:��J��{f����>	�)ĺ�r3B�!l�>���`{�HL��`���q��O�4B�	��2,�:�^����5�=�����;�ӎ�&�M](Jm�0�h�eF ����s��&T� ��~���J��p�c����iV�W ����7r$��_���u�B���r?��f����&�𡩠&����'fd�;������KR�ߴM_��g>g.fg�wT�  x� �Vq`c��xgq��M���Ǚ蒶�[����E:.Tݼ1,��{ޢ�=:�����m��o)�/	M5��p���qg%�?�����L]�m�9M^n �s����U1jޓ@06�M&�Ӎ��]Py���P3����ne��lE��O3��[�9/X.E%X�q�-�K<���������"H�0�{X���N��b�.��S�w0\��]�pz�x��l�"�m���t{��w%�͗=M�����?�ܩR��3L��1��ad1�0� BV��Î�{P�=1����,#���8ט����w�y ��N�NQ3�%b�h�p�e����M\4���(����'S�j�����{$�O��Ӓ�R����	3]�H��
2WM&��O_,�\S���1 ���p���՝�C�_�du~�6)6�*J
�d��s-�u��2��Tǃ�9��#�$����=����_�����ܝ��?�u�nM�ANcdt�ٛ$�)�� u��G��Ǣra�Z�K���Cß�����~l����j�w����\�M)eR���^إ=�@d2p��O=P���������i@umv�R�R9}�SN��