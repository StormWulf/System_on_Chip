XlxV64EB    282d     cc0�P�� �W���At�@Ŋ99���ӟBJj������|�9]~:V�����M�8;X�%��`Ƕ��t�"�8-����@�X;
s~�dyͷ�ʓ�c�������B'���{��x$��՜+�}��R�v��Vi�m�#�y{���!(��'lY(7������k�z�2���	�m� c
�x��o����\�O�_&�n�͈1A�n{�8[iw;�2���k�z��}x��PL��0u��y���h5l[,5��#�ac>[}4Ew�D�>w�H�[>ύ�=��-��PKUy�'�(\.�"Se4�O%b*����D��v*ĉ��Ku9�8�`���"]
�������� J>����\R�t�L����[Ê�����=�l���w6ɝ>2�������ˣ����r�~D$�1��bO�)3�w2J����V��t�ܘ��x��:ti����g�1M-"�r����@�뻓r�r7q�m�v���U>��>�NX8���p�T�Bq���緱�xn]�Ϡ�o���!�{4"��b�-��][x		�
L>*T�J�f�p����'$7A0B^�f�~G��̲io�%-s~��TѬeUo��-�j�^�s��q1��×(�l�^F�M~.~���)Jٰ�n��F�RM�P�~�/} �:� �"W����z$�,�����=�ܴ�v�S�c�S�� ����������!#I`"T�xf�b������C���驯���x��ܠA0|շ�R]�J�;ʃs6����NP$�%�_!ݭ���dMX�̈b�e�1�����s��W�l���Ʋ�,���3F�:�Bzіx-�|U�,5է161��4�b>��6�1�ڐ��
1���Z�t�q�0^Wy��l5R���T�,�Iw��C�>���'��8+U�&(��kĴ� pд���ѱ���E���9�����)��*�t��b
�����g��/oX���xŠc�݊��"o+'ȵ�8������P�e枌�O�d��&�[l�p�%�ϫ�I��.r}�R��f�`~��f���o9�*��H1nT�b��zY}��S,�����Օu�r��ƈ�.7�t�ݷ����m�q� �u�p_���ը�d��������������_��0�?n~�nt��F�Q!A�/�y]���a�����ۉ?���)�*r�Xb๧��jW��06R��fl��ު_��T.�����"���_е�:@�s&3H���Rr�lF���#z��S�L���wP�������mEO�#�k����R7�P�D�b#A=h��ت��3���*��g�m`�3��"��G��i��T싗��U�Osa��ɍ�;�@��p�%|�ΒD{��<��J��͗f��b>���@'�LxU_�ܯ<�H ����N��Cѡjˠ"�Gtv���"�rs�?��S�*�?7��� 9/`�ރY���9�Z6��ݣ�=��&V0Ak�ed�A��T���R��1y����6�6�"6����	Gz�+3bT�ҕӾ���Y�s� ��]���;D�z��G��&>?��Lnqm9�rS�Fu̖�U?*��1�~ĺ�+����UZ�.���В�� ��sG�|o]��BV2OEm+�Ga�vs}(`c�ݜs���i�dpu,Xۜ10����PK0�$)\o{$%tE0Kx���6	�ā�NPke �=��k����5���ϼʥ����7I���g�!CĠr$��tT���G�M��
7��a�V��_RV��L���(V|�y���q29�SY���mt�eQRlr�9G��?8�'ucԾ!�ʍ:���_�������eEJ=�F���N$��c�жzGV�$�T�����M��$�~�BD�>w�k�χ�m
�j�]�R�IW��'�5�k�^��Q.�/�^�$+r�va���=�"�6��Q?�Pn�0$���.�=Cp"*���b������@��W]1& �(D�b����XQ���_#��N��y�)p�B���<9ǝv%F����/$����/"tN[�ӳ$��1�q��*|���=��u�8�y[�����?8/S����@y���\�\����g�8����G�J�ؤQ��(&�#Q<�BjADl��Nv<5�#��4=�,�h8�p^gK�c�mI�oX�#��;���,Fi�t�V2J:(�o��ܘ
%�\�G�qW��XĪhy�5_�J��dn@e~��x��~<��OV\���j���ּ���5d_�j���{�=e]���V&���\�M�;�Y�w��S���&��=/��yED����cT���i��[Z}�	Jxw�o��\O 4O�O%����U��ŏ~&X���<�d >�1?���]n0+�޽��D3��z~m�A�w&8l���B]u/`T�����JU'\$��M��Y����&wk��*7�$7	�����8�C.Z{C�B���OTp}{�d��u��c���"�m��[�;Xw�t��Q�ʝ�wY�JS����mUWs�A��䒡-BC����(�ۻ)��s�=r>�w�]W�����Ja=�B������a�� .���1�(��^QH���x�D���J[+%�{����"�[����?5�1T��2�3�w��/*}��bS5��}[ீ:8�J�ą���Sr�D��;s��o�0��3Wb���DT���UVC�b^\��W�>Wa5 �����Y�"��i�$���o�s�PD�֘���`�����-�9$�à�Q)�e����^MS�$�̇��(G��A�I� }�H�!6����Y2HYڸ���X!���o���~B{��B��:E�pY�����$��L�kù��St�sn_R�@����J�@,Rʉ���s�MO� ��8�.��&�ч�<}�$u�ʬ��s�023���1���Hln?��wR
t`�F2��&��7|W�[�n|$?!���X=�1_��<�������_�&�D��%?<w�-T����/#$ڑuޤ�^������I�H�W⅗��ū����R���^p<�� ����q�j�[���r���ג�Π`�r������nI����V��Ѱ����}dC>�/1t�oTS��z��s�ݬ#��E��{O��k�8��'��ړ����"�Q�/8s���D����N�<����������$���i�j�z���z��O�.�ꌼq��;�sf��+[�-�SZ�