XlxV64EB    5d7c    1410[�Uu���p��\�d8�i����qDD��6�H+�0R��t�j�������-=d���ϕ�ݻc�)�E>��J�����x�bt���߲_SṄ����f��}7�bx76	�F���u��95jWr5yL��? xY���c79گsJ��l�D���ձ脻;erdF�(4�����(/h+� ��eg�������4)�)Q������&{�	P����e|=c��_�<-��DN�Ή�_�U��cV ;�k�`�����/ͳ�]�E֊����.�G|Sw��&����+��s���Q;g]/�(��g���/7V�N�7�hKȹe�Z�,�r�ŉ��"���v%�;/]菼n�DR�6��b�	AwIh���Î�d����y.$ @�����)f����W9۳d�ZP����!�H,�i� �R�s���l����L����{m��ۭ�}��R��$hɒD�-f 8�M���0�l�)�Z��ĝ�U N�7-O�]ǰ�&�y�\�tC��H�)�<���	^�����9+��*}�޺�-۵�^ufJ���+h�X�6��I�qP%5.�K�;���#��{J;;UBrZ�f��f�Rt�D�PPi͈�n�Aʔ@Y?t���B��<���v��6���,�h�j�v�t�C�3�.f��~�)oQ�2A�`�д�T�JAO��&�{�*I�E"p��AO��uZ�o(�c�<2��2U����bk���`?B������{9N
H��Ħ�)�c?�|Et6���	�����@��V����Y���s� AC�H^E Y�v>��+��L��Lox�i��d_Đ����=^k]]�G�m�Nƍ����c�T�7ޱ)��:zМ���Z�8�53�P��e1.���p�C#�i�0爥b��X���m����~�[)H��\����[+�s0�����أ���]�&�{�ƿ��/�Y�-����� ���i��g�ܗ�{9aܕ=��tKu�c�]��?/::e��~��lkw��c�����ml|m�IU�9a��h���#<%R��)Xy��aFo�;w�����Ŕ�Oh�66q����Bg����(r/���|C�zY���"v� �q��Yf����*h�d��<Ҧ`-aȷ��4��Ռ��u���S�I>���#�����y��/�%S�����2z6�G�Tw��g>і�E���t���ֺ��b�fy�t��Ƽ����M��ʜs���<W��ʅ��O�@3c�$�2c�#$/�>�C����,�#�Q"��R��^�3_�S��bvP^����A��5������}Q��@�O�� ���G��C�~�^��G��A8��ǽ��vj�[�O\�Ԭ��[�DX�ذˤɾouʻ��X�[s,%�Y�����҇&<"ܡ�|�;�2n˲�W�@�5 �)G���&ڊ_l��YGs=�*�f�
p�đI�}���g��5���*C|���=C�Z���z)6��%��4=Ɇ�qR���20�R��%�0�ִo�/�0$g�E8�
�`v)�zu��7 �D��� �2�ʸ���2��ӍU�t�,��)Gn��Z���W��po~�$�:�r���^��*��Z���|����	�(y8X/�� �mD��{"���ş�N&?���GD$ߙdZ�����Z����1q4�ϗQ���&p���*��{}�}�I�c7�b�+G��Zk'/��h���9�8
m�0��j˗��iP��%���7@�ŭ!�g�0��d�}/��[k��W��K�<��ΉT��q�R�_=�F2.��M�2w[���E �η��H`�h�jK��Jeӊ�)���Le�����QN�e,�6&:�R9)ũf��OGG����c��v�zΜQ����3q1E��n�������d���75=i��ߋ��;Y\�ڟ����:�0����V�,j���C�c������`d^��V���r9=Dft�r�DO� ���
�2K��\@
�kJ�A)�Y������<�\@�@*�+yv��|v"�=�t�k=��!�}I�O�c3�K��A�2�{�Ծ�O+u�Lp��e�#l]Y\�z�r�aX�Kr�D5�a�}��zz�1r���	�� �%�Ok��z�#)19�KF��ئ�48<0ϟ'"�@ڂ"��񱝳{b*��ML��b#�.�ćą��7$�.�/U���g�A�̩�X@t(�x�҇S���+��
�:(�c�K���~\3K+NIO�CM�.Wfn[%���+�ki�
�[t�lH����W�`�Q��ř���=���!E��9�/(��%��2�j�%���+\�:_��`!+"���`���S��k� `�M����7ZP�l>��O~�um�5pe�|���#����#T�[��^TV�}$�����<�\�	6y�]�x�$�MfZ/7�cx��hFU]ME�dsg�~��B� %߻,gw��eT�Wc��ٔ4!�|�L?��C9���n���6e�<&sl�v}��tց��@x+�|�0.D-���������`5C�hm>�C6t'�{Ҕ�v�
+/w蟭�����"ص�����M|��̋^�1,��JϚ���	t^9?�Pb��f�*Nb�@�r��v�k��;b&���v`
n��&3�Q8�&�x�R	�J����l����D�d�O����:� ��][��/���~�<�M)bo�OW�m�V�����:#[[�#�\0�.��~���f D�f�v��k����{��I��~*v����X%�!c#��=��L��T�+n �'��t�����kՁ~�R,M��S��eDAj9��䗩�+eݷq�����+�A6X_�3��� ��\���G �y]���1jq���U��5�z�I�"S�o��6 ��5�e~>zp�������z{�%��B���mm�~yD���FR���i������6�	ь��Z����r���$x��5X�D� S\�5lK��gLv4H�jc!M9�%�B�h)��wt��/�R���f�1�p� 4��L�L�`F��şu���ħ�P�@�#��AP����I��Ylǌ	�<��V`^-�S	]7���JY�����M��^2R��1�s��Y��Qf����&���4�ga>L�7��a��3����?�ޖ�H���K��	 4�p������\��~�u/����p[�F�ʞ�����ۅY}ڼ��~��,mw��b��l�	4���Yk��[L&��V�X�ա�����1yG��w��3�*�x���va�G��p�����sF0X��c��I��WM�Mk)V�W�<(�������i這]Ѝ1�->t8$���q\���OD��>6C�d��p-�)|{��Y4ɿ�E�U�w5K_��l��������_r��Z�R���E=k9\}߷vDӝ�>H>��mȓ>1O��%�1ա��?�����T�YL�mw�5u_��6�����CX���J��W�ߕV%0�np �Z�0eY��>��U]�6aÔ���,�a �h�i!ȢPN��^��2�� ���d�^:�ڸJ>+�뭍��2���L����H��VD�f��N�{*حvJe�-S��(K� �b_����pZ,�}�{Q*|c��$�O�Y2��o�&�"�[����}28L�VʦN�O��:]��O8KĀ�dЩ�C`�[ʭ�t��R	b��}��q�-�Bʦ�O��h�T]����W�ʇ�z���%}��W�t3�*�uB��F��Ё*Y�t9�=F��W�Շ�m���ȼ=ǽ~��}C�kr]ro;&���%�W�����g9d+��$�Lgm�[�����9�S�@?�Gn:"Us����WB�u�c]9-�d�.��3ߨ���q�|Y���j ����Ժ$�acֳg�g��Y�)"y���GM:�MV�_��]�M���H��]�W��ա&��m�e�ȼ�O
9i�=*bf�g�����6Y�!t�����ci�nNɆ�1��+��nn����\����L&�l�Cs
�ɩ��s\�<홷��0��
0/�-��a���.!F�xɝe(V�OP�<#L^��iK݌.~6���_~������.Ӎ_����=ƱA��}`
u�1dֆͰnaF��]t��,^����Q#L�X�囈��		(��;�p��>�>�Nw���Y�������-.p��} A�bC�c���M|����i������X"�w��L�_����k׍a�G�4nHANA��q�5{b�5v���Xx�f;�S ���.6���D�9���j������zp�"-�2�6U�3p�$�|ϙ�%�C��dMP�d�Q�ݞ�Q|���7�%�L�eųe}��CԇL�љKR�}(��4�����|�����|��;���ĦE��v[����)��z�R�G�{�d��"�$�����f�Ѻ���3�p�Y���Qo�x<�^^-����Ϝ��GӑY���T�3�Z+�x1���Ni�p��UPd�{ڷ��G?�G�I�N;���0�� t!A�M��M~��R4U��S��g!�����=m�Q5��HIC�DLI�>\�k�@��\�ג�����=�hK�zXSs���3k�q:�λG|��W�	�z�.�ξNPlC�fJMH�t�:�B�
W~|��*"�&��ӯ�)�E�I[`��Vs���dE��#ˬ��"� -�}�_"���G ��W�e)��-	d�i��MD�<㔉T��JW1M�Po�ecmWd�5�)��QVy�x:��������XN�p;�+$#,��8d�4��Mކw�k�{5{��&L���;=e��W+��m���7z��rd���y?Dp�-zɳV`���_�Dg��������.n�s�Q��aٞȨ���7�D����6���"e�уO�1�Y"�*`���l��|��U`��
_ڽP6��\���4q��������zmU�U9U}��?�2��^9��C���.Q��?�w�4o�3�Y�Q=ow�]|`����4